//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TFvPjZP5fpCkxPNDwLBnny+vB6d83sFSsyL/hyKOIXgierX2DQJc+Bv+Tr4k
8KPhWya+WbarZXaCl8ZzOpZGyjGNHFErA2+QiIyBR4M7iwigYrzIGGQqz1uW
ugu1oKidx7jQf49xggJr3SYSguuUT8p/p768RjYjWPZEo8z2QmqkiETxfUg3
n+1TmkpquTf65adWpjCwj7EWAoQaZADLR+KTgFmE3BJ5aEknIIxc8iQPNerE
ZEHHMdSLDYCZ+N2cn1LEfSHuLI22TYwbMQEZpX23Ogdw2iRHxYt5xjHkC6rZ
9ug+Y6Zz9O32wlWYyHXmUAHNm/RyNAct7eOHVDRcKg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MgJbq6XowQX65kZ3N4BBXmQZ+v0xsyhPfEKviIRaSwHT2FQ5T3wtM3bPsfyn
7L+7agDgQiJxOx3H9jcOCfU2y9V69xejhI6kKZGHApajW4JOwVLKDC7L1FsV
I1u1UfXWdxoRxR5q0jBaEVNFLdXjq5DhpYlJgOkRntGT6/5h7IrJcoCDopuF
z5D/WS+XFxnJNvcNglKLfM7Fl8KE5nwm8X4WB9MDJtCaTP+6N1D1KSUXONy/
CzXLO8MOI+1AbLF84oNr0ID2bJrFLeWTgX42u568QzleuSUqDk1gN5yTRRZP
diprV4HyFqBbsQvb75l23LqqC2wtDSU92lgzKS6nlw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YgeNteCqezaXje7wo9+8s2u6Twct9gzMBFdBp9IkOFbQOZYp1MHtY437SrEC
mi240rIwyoNKXhS2A9RCRzehok2C8RVv9V2ptuYk1hAhJOnCvYyA3GGukEYt
46EGPrGoxFhu5yTZDmFh4kZv4qhLyDm6A71a/gSZHdzatPifb1JisRLKVjjk
ZpS5ArP5EUBYe6K1KjvZ3hJOR+tu53LcADYXrVPkStbh6Xa/xVFe/fusKE32
pK/vXkq6DOG1yErIBW6XBO98FXkByHCew5oj1077HekWzLMdZPqabyM7U+PG
CN/xUNQTsD38MOB64My7utnjN/z86fnu4RyQYoykyQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NqSyJPg+aNsC+nkG7gJUO1m/hRh1kWFpyVUEJqQSF8VxeXRVi764yOL97w/W
bGEFrDquVyJeSXbxzQMQBoTCHWcV3/P43q3HfU5wRZS1v8p7XoXnaxf7KTBX
Cec9jnd4YYAdRwWg/klSQHKDsI5ToiHndaP7HKJCF0oBPRkCr8EQ/UOfWV5V
ikzaW3vqi7QM6Crwb6aOdx8vmgsCGZsfrEgoPRRfkfHiyG4EZ6GR1XqMoIfi
7MdMlG4kqhv8EDIdSDXWH6UL1FbdfbvYUElWolujzOl5RcIco1LNteSv0gsw
tTDlQLmO4eEkWgP2lNc7Yh6YonkJ6tyDyysTFPUTbA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I5OcpRAhKIleAsaMju9jlEaQOcUtjVTB7tf5VXum4j86mBwL8Gh4ltQySZtW
/DvwNfIgFxCvBBTJzgSUneECSgVTT4nebrpBN5F3zAivLXgMBbn7fLNFuoWG
VJDVavc2SjL9C0pGDP9Id4dkYP8JrUTC6w0oYkNcskxfYwH0Oj0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bLSUoVfDIEBkqQduTlOf/EYxSzlW3I6fy6b0sf287Q7Os0TUeM/0WuT0iW44
hCnsREzNhTRUWkvx0bWZTULU26z2yg+W8FwfKsP0rBtci8SOf8QXEYWPw6wU
0qL011lzx2Jko9epEu5GF1z9iYseKTeNqialcZJ/87+7hf+a6pJEnkRpG1Sx
VZIlUuayi+UTp4t65b0ZoPLj9ecBebqgMBwKIGeJ51YqynmEEOTZCEq5v3IO
vM4koOCAUq57bVRWpq6GDDH/8qnfaKoRxQski4CehBkyX0jgqXcfyuUXSJTU
jxTl6WrzFxiYtLBCAUV/xvA1bzzGiG6uZpo2JAUUUCSdFinfmbs4Mi2enAaO
EL97eU6PvzEprzdy1MvdLhdegxHD2N+sXeQBnZ0X8RXb0k2mCOJO3yV9A7U0
Gc5fq58KI+mn5ZaCwn0fdsNlIta7qeahgFCCz5GD5oBhl7Lq/jaImnzRymUw
EFQ40xqYF4x9WFXuRFWb4baxXxjey6xk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XKoRqyACgExa8McY3yCTdCX4MgXftnlT1TAXNPwk95T7OMmrohn8mSd2FtYg
A3wWhVcUz+wFCCuFYwsETVy4AQn1EhaWdV7Axl27Ewaejz5f8K7Fg5Ar323a
2+8DGxUuxcavbeGItPkWpfqM5RK+n/Jd0lh66JLkxRQwfm5khtA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ay0tvi58SNxdvnW6y+fhLOqaRY4u6IHw81iThQXmc77pHJhUGWnsGmIU+IQD
woTnzCOb9MnYGvyEtLIONFEdMMIPqzXykTHlVsUdg/7Sva0Kt+YHrVtIxn8x
M9WAWEpxGBsO0lW92LqHHYlv18M1KZ1m67xGF3sgDXG4xUFBXM4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4592)
`pragma protect data_block
CkJkVKaT/5mLBM6rMUbvzKED2PQzgEFJSv6RZRgc/ukHxZnwmqkl5kuIhBfG
uexmPb23216M4h+qu4+kTXTCQiTq8oIa45f5pUgyd4DrOXvwGeqh8CegkHI9
DcMZ3y79oYs51D/fH58u+/dwvJugJVI0wvzxpRPS9Bgn/SIv2Rzg0CxKlV+O
V6rNt7b+xiCfx/xJ71dudnURqbDZEBBRjd1KctKRihRKYyNAF+XxN5lBHmeB
xxSwGFIdC3jIfzjKH6AXc8lvaJseL5eIhqOGPRsAL6KpxQOED/dkUMulpgZo
OQ3FdvBg2GLo0aqa/yetQH7dOUXJLu6ML0iH15M7RsSb/1br9vbefYK65iRz
bJByBlEYSpMPJRNXbC9WUPCS8DY05AWRx8NuZHsbl9tP5CgQBkmxPlVbjHFz
xniWuazR5qGwWP3V6+sDaXwLjbJud4TfUa/ACtjL/NNVybHisw+rZUKPgXx3
L+SMfIKTTE+xAZyQi2lbDDErV9OpW3lusyxjCjhSa5RgxyZ9VsRXzjCHbqct
QNqg9IfnlzdTvoTH34tqIxWiJK+2EAwuoaHf2ede37g2P25H+L2dDBZr5HZG
EQorw2jRPukY+lPm6QlthnvF+mPkeMz4RxLAm2P6IZiXcRe3/AgnmkapwBUS
g7yXtAo9xsJPIhVY+RwMECcS1zsZpMIcE6DBoB599HCRuFybd926H2mQx6uL
6jEF9WccVBqfz6WDXAQQR4PKQEvATl8sVT9NK7wx6xZpejvQ3K7y0MSz/P9J
zn4VuG7/1TCFudB0HEvUR0o4z2NNlO5xC/Ke20Hcw60ng4jJYOEp86LzcODo
WSrqPV0n9oKF/PH/pjHHjchOyqg2fJWLKSFmVEnLZLYs3jJ4pJSaNAI2nEvQ
Em0JkkC6GTvKCTCoJyt3Q3kMmDGsQsaBbC1Ha3p46wnd2CWdu5QihfE2q2wr
7BKaMt6o1Ll2Ks5b9ZhlhXMijhBelKMTt/tkMx/FJlnk+tT5Vq5tBlbK15LC
LIPrep9F/BDDieUX571gfpqustzBIHDsur1blt2LYpJtmKegFUh4eITinWek
RFcjlnMs9w5Jn76LxDA8LHk5x7kO431ZDwM3drH3h7hxkFJW3eXoOo7pBjMt
CAEm25ZBQMchsS9QMMTMwYGi4Rj+pC0ak14WbUyq6uGGlHyOjgKzXBeme/8Q
Lk4V/w78UC0E+91+ddE4hkPh4nU/CWMsUglObQXnMSMrwhSj9KpBsZbfAWxH
zBroq9yPJp0RxW4jrsngzJUUheLq56A2mPeCLCY1TrY1k4uYGvMbMwYdYnXY
MOZIBz1eUAUoi/o6UngyqR7n5UtegJUe3oL5MRr+4P76QmBX4UhKD6Qjpn/e
KxG6gjgnLsPmmIZBmd/3WqB9wia365cLx8ZYb69X6ZMivGF9YdmrVf3XumLj
TkM5QYWRobnwMOZa1F31gjmBqAFshUfdEXjnowzV8z6Y704F75z6TdULiz0+
EgRn9fRvfb140HjRXJludDLKGHJ21eWB4kS8l/98BC1Xec4PAYBKRrYVvP5W
JcflWU3GzWC8o37aZPuKYkrZTHPSiQoDkBGh7+nlMdEPlV3/Ugu2WxRLUbLT
kuecMZLOcl+nyuz57spyAEQnAv83hGQHVBbFvlM0FIpVuNjTeK369Sk0v8m8
wBY/l33WhNFscMu1XkQ1HFesOOUwizUaKyD5KNLo5FA6ChUuGkBAPBOxMNoa
CAxY0SvSED1mtrfVI3oUAuTXpjfmZ4ME7QH8Dy7cGLZDT4WYMFMGFJT2niFW
4AlxFmhMjC8ogMVX40sXLPlKQANWFOw9WVJz4KAv0wMGGLS9huV31mONsCA/
ZZTRe14eNRUCwjtSrsua6q98YQjNlEoGeiz83NH+EfF0iNtOPTlylu3O0XFx
CzEoRUPYKCQpjFhr3xdQjo0TIj0/v30IVDmdKyLYU4y7V1OPglXBCRJSGjjL
XcGEk2g3b6EqgU4GznNjnImo2s8LHUfQhqmLBL6M6N2PwrM1yUk/oUxygMFI
jVttruz0+w12OxjzOq3KtRxfjgfyz8Y/36gIF6bsg9SwJwrDAOHWay9AcLqh
LeJWT2d7UZ3m6p+JJ+eyQNX+MVo3SL01QOuEhesDm3Q9DLLVR49K1doKUwo1
dlFRzRIiDMt1y0mjL/QFZysQDSdFdKgyyYo2ffVOZPBiHTsMGvLcxOOepHAK
oniEO7DxZKjVgYtM6cNJpjec6i8T7vFLhU8VjwWwS1J/hSOLa43uhvR6zeRA
p/dDqk3qIt7nb3fmGDEnnOzFiaAhpHyRlQBy6jVTH6lDf1qgbZZQT0Abn/Cp
ct70vf2yJYOLtKWkgiKLfgLL88LebUnORhiWB9djpYranu23oxk4r9yYCPRj
jMxYHleAGwnrbDmKCbWbRJ/E0gC3fWXVHizbcH6g3m54B+IWm/CYPwtkQ5QJ
9iYCHd0Ap9Dubjmsz6mt/T2uvxiUysJAW2oXLmZvlpJNhS7n1wUl9QnqYVKu
x5Gl4KUTx/PCOPQjcEJrfkWl8oPL0wi/q+OoPmZitoFVpp3C+9rWEcSYm0i7
+k71WnAuL9af74TcH2eC5SIgCWGcJW75e+t4aA4wtQBuZy/H1gcR6i0ugJmi
Z43/EYjADWlfn0SUkB3xZDSnrlQt8A0IQcl5hcL+OlKGjl9KNVCfp8BxMBA0
Dzwtr7km4aooPlWP3BL1dtrcw2y4tRvS+38mbFK5Fr65OygTFyEiVE+A+AdS
j5jBNPoA35TZnu0EqCp/AXFy5aVHTIK1fvm2ELXuYN7133J4nrP+M4yWzAdm
vw3Gz7NW1JZDgnVea0MWROLUpko8m3472pJoHlT2YvvmXmVu9DA2/bA2nyUM
6HmqIgkMT1Ea8jWBhc4aR+m4u6+ACgerMoITAkvVyG8Z4PwdZG0m05NyUsdN
i8xwkWaUoIB8FGxTuJFNMbpT5TaaU7ir1yVrHmrGv6IKyfHIzCKfxYdvHkY1
MKn3daM0LeEgGBhXgab+CSDQze5xwugIEghxjfHkDF+qD+bZftAHYEbOpjk8
uOFabk9GYMF62kuvyEAsRfQDxR54gDTzPUXsk79mFSr5+9MJ8uyF29v/TJls
qmgZQDtZf/fSkexNoH1bWadjIqriAJhVK37vVMHurFKnB+ffSgfXpQSL+rx5
mGkwDPdrLagthqtpVx0exmyJDNFlfON4giKt1VUHpCvLdBAtvGmaHGf++Qtp
ZgNfqZGjWe5eZr8hK/S1DuEz00iz677ZdjRPXIeKKXcTpeaPncuj9+06R6rE
AvGYwzXK5RkSYvyvw/pmYI7G0SqkuPUej9OdjchuKY3CeflMe9xEGsAHF3yR
UiaKYDuA4DikOTI0YTIn/ctqlg1gUL46LUb3GMo+RSqiC057omfn1Wez1Yte
3FgWL+aBypAGC0w7w5HIkfONBemDEGGcmUDAfuDCFhh3gJah74nxeiOE2hFz
HRS6HZds5/zumvup/ECtPgscKYsljHdNSkZgqECncqRkzKsolC1MyQ+TRJyP
PTh4Sd1i+MFzttoF4T5LTfSPrQz1CVqLKd6lzSf4ggxQnzvH48yS9J7B8tCT
/JWHkoUnWALarbJn3+vGF5PDzN+HECiMTY3ipCKDjvhyXB2jiB6v7reeVHms
4+Ydku+y+NrYC9kZ6S36X/R6zGTJRuTGxbI+8AyH0K+QpyCVPClaLwVpsqdi
RpFMQbVGZA/qT78t7F0B61Fo9M7EgZog1iZZEvAA78bSkVjneIj1YhjxSC/h
9mV76K2sX+WrdfnahkxwE1/yUNcRsRmkZxqk5cGDQ+6wZIjuH1DDF80LivLX
Qpeamv1MnrMYbHGAPw9zI9tVe16DTAUf/7yKC5ct/UTMaDaHJaMs3zlY73J1
rGIqSkdU4FDd98lHEbigEGKlmnRZZWHrI0+aEXpWE2xQGI5DovzSJdq2QgbP
/lL6tmfdsG5V318s25qJ388PtwA9Kp609pDCG6nROlMnRvRFEjdwvWkYiJfF
DvZMTDetqiV7qHCJgjBuq61oqSOjVEhJoSFKmAfwB6spTAFUj1A9bPGOF/vf
LRtFX/TG3jUS05E/O9pLAs9uIHFQkfj8M/K3P9jcf8IMgsPO1BosyYXFVW/+
FtFSTP0sbtB8xTltllRNjBKRr/8BQg++4zfUaz63xUWxe1438f1omuBuXhp7
3nJhtn501shbQuYPIPHfmmUWzdYLbGl7gpNiSg1t9u50PtRkUuPy1X9ywN+S
e09ggtUlUPlLAyaK2klZiTXbTikpBgkgmBn+ZX0kAu2ffbb/rqHAWkyX7ZmT
MjElJilo9Jb9f6B4sq4chbJ/R8AT3OuKIAVf6M/ARFdWA/rUodVoF5SGySTn
O45tDv/1qbmhU5bovqZAiOvZlbMmSkqjPsNLcEIyAWgIA8uvd9GxTubZ2hz8
auacL7srbaqiF9o5UBlUV9w4+GEbl3SOMudqR9u93O+PpWnXy+LvkakE9cdA
TIQWXaS3DASnrm7MOLXULQYyGd6fkADs60u+FKfl3EJKEb86dguzH71tMJoX
WynRq3USAzpLdo0AJOnyFUwwgj8L3xKt1Wmva+tZ9mOQCGmJIDDiuLxj5t20
w+XlZBBlMc9B84GgS1FoS3yPs/j5g0Zm+iCTM66XtZzTUH8pe9Z3OBgGtZuT
dHTxECZA2vwXIf8B2i1JveF3cpG2DUmjc4pz+ddY+Q5f/DJIlhSLsUVYF1jI
uJtJvaSEXcEQDUUIwWPfHxRzpYjdV4x6x4nPQInj/HBGLYZFw6Spc9UwNH3e
s4wTPhHJgb9Blmxp3+v9HJ1MShtgqcSn3oogr87trLpUUDxg6SnhMu+n0+GS
SML2i5Ew+t3A/3mgReJKhLon5Ktucb6SOHxaqR/wuXZIQHEMefr5/fYCkZe4
o5PLIbsbrCWubB4aPVJQQIFeoRSUq/oBV6nOEy/hbLpNVZkwg/2QZQT2wCxa
WFkRYXyyK1sJYawNk/sLNfVmzZGbCK4kk/5AvCkvt0ICljz6nD9bdhf4A2XO
NU9Of9uKd/D08YM907Xyzctr2MPUBsxd6e0cebjzx/Y6rPBrb6Kc0HkRNvJ2
EtCsu0aBwLAuMlqK36mxB9BCpko795WewVOiZVNXYL9Yqb+sZeEpZwK7BeU5
2ppFK3NSzuPdSYm21BtjNjLJlENEG1rnsyA2Keci/woRsofim00o7wQC1qaa
U3GtygLhqjajXwuYpf4qNXzoIMkvpuBaowOd4uarWrSnIKvClOLB57iZaMzK
VDmYuu5ThmwncnPXUtaOT7cGw2paZzh1dSLhnP3twYBN+s5I7hBIGG4dAu5w
LeULVbIT6N8uVHIBU2dnpQujiHQtBgaEQ2+EgPoW7Jb+CbGkIu4FD3AYtpCT
EXvpx2K0MgQiTO4tv1CQ1+o0CfsEw+SPLTYim6V00IE3e3LtLRR6wmTcFnwc
aqORDg57DX/JnD6EuOYPEqOP0uJGNCl8De4hJpmN30z57oE6dxthvQE/cUOh
eqruDLutJywV3ynIEKNB1/PzDXPbVleituYfW1nMjEOa2aOPYLlpwoQhcRVn
K28k7t1spDhJifoFRxBQUKImM2NnRiwfPg9Eo11DmI5UUz5JHsLlR2c+k++k
4dUc/N5y8mHIXzKM6cVfAngddD24Qa+ESbX3wZAlK9z9a6V0Pjmz4afRe23j
wlOyPLB8ndDpPGGzQi2Y21HlPYAmyePe+ug8opkWuZSKbp6o8QZ/VeBnPhKB
aua7tooWgsTZ/fGmbmph5RHfDG4Li5vj784gLed1Q8ZCvm+Xw10FR9n8dQj/
m8G8MmwR08DYrAST8xH+V3rVRu0YjBLPjIqRehiXYandRrp9Pw9okoJB8C/t
JvFbyJF1IFjpk2PiFZWi2C7bI1217m0T8csyuo46ELTkPq1vpVC2HpdVIbXr
qogmlOFt47aB8cl8kuSNZquAm/LYDqB5NlAPazsAa61RXFPbQFvtg8zWFO4h
MKrhZ4xnKUGcDDZkHmri0NFoJjefsWbrCgjYLoiJWt7Vc7qMpRsLFJ7C9zD1
8QF+QPpAcRCG+kbS+ea6stQxtlsWQJdK7QtF/i2jgXWJ6ReuwcsLnvomcgPr
0uM=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI3Msc29mD4DEdaOX7T0x00v1a6CKzFBS8qhTnDce8zGrpSe/FRLTSTvQ627SW9l1bK/qd06ppIHdXcoxJiZTaGPQE8zOWB8MX+xVdocLt3P5PeAlm2nBnihlneoQlVp95PjJa5CD4nPYA9nnW9N13cQtW0rVJhZm9hLVlk/cTL5m3HlRVxcGlNiGD6/6spX1v2BX1Ytec7xZS3MUVkooFbOoQGtJWtX2CMAJS1+K7G5k2TCVk7DRmX7aUo08mmzxIFlVPtMxXeNRgmjOGwmyQ1DEBAf6XUK6S0XhBkieeFr0nricH67hlUIxsA5qLJqI6r6HK/2yeDzrZbHlgXLA02uyUQ0KZLkcIULij9MLL5txH+EIAPS1A0DPOA5YUpWDlE39xvhqTru6C2kQE8hVQsO3reZMurLIrNzVzz9uBNmsvkdmWntsDQC61OBDHc4FOU8HcR7qL01z6bcEKaQTNQljIccwj351u8uY5zi6RxkvCy+BUi/obMchU8yC1o5yxrOghmTkhBdU1vwEasPLyRdrRzJO+myH0eiOuHNFDjQTj0IdXHlnGRAphzC1Uk3UdfOjfzHqBVgGLWrvqe5vlrmvW+dohgx5gFo0U24ahaptItSxJtAuwGxvVp1Q3zZG8k1gchAwGQ/vjKzoZou98MZlAYlOFxjiCNX0b7MCaPpAyW7KkbEpl+eiVeBJMf6E2kGTseQxvzdX68nNGYvKJx7JSzQ7z18fwudHrsFxCJq7zfbz7RRmFGgovJD3r8E6kDlcG3hOJP5vR+I3VTcm4pv"
`endif
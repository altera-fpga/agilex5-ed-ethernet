//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l2tkCFccUsRy0uXAnm3/EKhn8AGKC6nMKvnlKZZM059LbKnbqS7qWIszBZ5N
Ia9E5T+gVgDT/fe+/2w195eqV93rFJL73pdOmSk32A+Zo7S9kja56CXdceUw
N+MnAYbgZRn8X/OBOiCBgOD20dfhIxbNnYbD9dLkIvQ5xcABx9/EarWMaxBU
I1+zZL9GhyRAk0LEY+rfSJPrHNlqVWngnuJwoHG2Vrs8nOBEpPoZpVOutihL
YyiknYSZFrjobaujJ73y06hzbPLDXd3uR1/zjuLHRGyD5qJHQaQiuvZAfeou
v/VHDkAc0eUwUjVBNPvD2oIwdCCWjKrIvLSEhwS3tw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lEQyY9RHOZ0rFTQPIviE2tC18qZ8/4Rbdhg0+8ked7/mqnPomK12Mfe5lL/F
KdcprD2cSB5siHSnWhVnqjjAZx+UGJuaD9IXqkRnlHwAhBT1/FdNuVuSicbn
+cFcJTf1rRuSfa4cWUYSwxTITq4HTs5Knz85wRA6He/ZwFM7Y7xvWnLS60sj
oBaFm6+d7ofAAUfFxLjZl+sbZA2spSv5FXlICmr1851xmirdYUtWOrDbbjAn
iuEBvvW0XB3SX5OTDMpTUdTgyeYWZ8yYLHMhxD64218LAkawMlxHKhYJW8td
yjZaNKovZv1Hy/qWuSUZ54wZfprRM3XpQbY/5m0noA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
huuqDkU+lrgMRBoV1opoi4jvwB84fpPtkeIKw7jdxgJIoT4xNL/jpasIawtq
vgAn4fQzgwOD9fbOuuSQZVSz33IXiS47srU/53LcbtSZ99UMEoeuz6qKMBj9
LDlJB5MDkBASzNo4bJKE+flVVme6NXl6igXsXluNdicW2yeV1SkULg7pdKt4
ww5COyYym66rxwpy9dFV+UOXYolx/vMwJzTqpQqY6Dm3g0Otm0oxOnennVDb
Hwzd+yZnTxZg0UHvshVC8V4D5yqtyjMJc8U3O+w1qGnv425VHS1VCsK7FnZy
ZEqaPSlzesYtB8KKjP4ffx+6SxE1LzE/5WOea9lxOQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OJw9Z4bVQjTaaSVdYLr0kNLhp1TgTxVu0rlSlebRo3mJ6CPXXi95sj77ag6T
MO5X9TNWWGHpi5jvA0Bd/KPw30mAgRCCMbBwp7aCFDiYOSTJgoCsR0AGByBc
DiXVdIcrsDh3fWfRwZkfFX1oOiIgtWq4pAPZDfXtA537OIs2qleO4LohiaeA
aLKaLsV4Ez4Vd/i6c/obgWeEvxMOeWvkrPGZ22bH5pb687Lenk8SuJd8lX9O
LMOuzasJef4Eor5XKdf17cc5idOHWCXpQNWFfPwNuh/5tXYkcZ4tyHTfQ2Ed
LQRep662TZhbV4Af1OCnTQfgicYInZUX2tHdEgCeNg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LLxbM4YwqiL38SZC4+oIHLqqv4MK6mdhl1TUpEhFdvPdN7VE57gUnkcSCWlD
WUSJaFVGHG5yVHxC2V7LsqVV4mR00xOD74mQFI5ELmjdpRN22e5KHikI4EVO
Eb8fuLq1L6b9XRotrMH7mkX5LHbDLAgJnhOxpQS63kJzOdXhvkg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jsfHw31HDVJ/WJgXMhNOFZljMZo8I6XbPrdTmgT8hyUx0pRBvzjiX/z4hLzN
ZKaEn9lJjcgMCDaOGU/DNMI83ncEYG3oz0RNRG3y9Q91e8A8S6z8+Xw3/fZB
Txs3iyoix37ZTWvSdNAUfeUas5IGpJya1fOR/X3/NGlZclPnW0nP0ObXvpY1
b0bjx/gohv2cY6xHAkBUxRJIlZh1e7Do5OYzUia4XY/HAdnu0sDKHPRnH5qH
Xx2nHDNSttqAgerS6owgrTinsaAY/pDxCMqVNNn5enLEMt9u0LQ2kZ5oOktH
NBVLzRDT1hrDbNVf479iGATBKh4DAQ8yJD1N0hxWJXEB7i0BQVNwwyXCf8E/
XRK6v41QJ+1lX0KedbNKzzbBujGroKEdHZ6eFKYE+a6c/kY7CCt1Si+nwjV4
9g/GtNYBpEFUeJmCrMiQQc4c3dQALKq05/GmvDYRBeb3sO9hp0vRsZixlPZL
2V5J70Ae2Dpq1QqbTWy+MsEx/IBVIqNw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
imtlneWamDMr+LzCs/uKwPeyD0QII1Ea1tnXKvIL6hrBAQNohUMm/GErilW5
hSblcqX2TzP1WX3o0rxyHVQkMV3fIWA1m7Dkdc/oXk1KjMrUcxcC1muZKSaI
AUh7aRgXMGktCWwgpkyp04lbGoXLG58383OTePudpPCttticFiQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L0ZKNpga+JsVhnQ3QrJGAx8+c7tFV1YLljv5lBnvjYCmSIz82QqhuMjIm35Z
Zm8HDREY3wDB8+eAeWVD0lx0zSDEPEtaNYlzuFi48RE9PgCJRyiUXllp78KY
S5iJ5NZXGVucios0kHx11XHJgsHofSANf6ifVkRu2TAOy3R/lYo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7088)
`pragma protect data_block
60l9JRAE0BAQoCu8W5nKRUah7Rzg4GBlE7pHC9R5UmXMZXadkv8/lOpOdNZJ
Kn/bIvKeeotbXTW0zKWdQbPyQmydz8rX5q+Qxh+txVY8epwakhNpIWYINtm6
tFkflfJHKAAOdXQFQal3tW3i1slpgsW9hS06chLt5ZFBA6Ugwvmbvp+pyd/6
0jLvcITL6a6HrUb+AjoLHWJNl286RSSVdESofa2qeMVxzu91oLbMPITwJAuc
e9+1ZEAuJVtEfn/U1GoNZ40JwPTRzkYJRCklVnBf8Roh63ZZ9nM10p/PGTQy
01qjkHdPhOt8lrIffSDSSP5WrRdK1vMqgj5+I1gu4oRWmBxSGr9mWwMEbP+7
diNO4S5iyOYW041I8SSU0KPRKNWGPttHowmu0K9sulhBK+m6g0UlIHNQX0WF
u6BRUG4F0+B9Xk99R1+AIHp3J66G/u1Yfy1AurecIxb8cSNUyV/XIjuE0cXM
Ef1eo4x19QuO5zsgOz4mHQQ4cRlUw7ACIeUqH1D9iOh6B0wV2k4el5Zi83G9
4rS2OpSdoWaxYqETi9QGoT2mfjBYpVVv/JdRx6aZLC2RgSoD4Z3op5UA+xAe
9/xLpq17QTrLvOHqpqanTz01IfwXVtMhpH9SvXMFj+kIpxgar/rGljiujrkO
KDb0E4tjQidlws7qjyURrI+P3atIiu72ZiR+qtyJiicc5JUDMwP7pXIg8XUp
j5jJ+MpGY/nKEiaHZkxW/Rb04U+Z9/7V/X6HGFE4UoGnZutCjkeUTpwi1mWv
DcT4mv2zCZG1zvobdWftYuqeRTcsr1XSgUZzsfT10uNB405DydzIuXBsMhyP
3t4EqH8iDPtSI91tn28nbrFSCROmr5A4DBGI/KXmVATVxi+ClSoYzgdjQfrB
rzW6RqvFJOr6Mr/S5DBoJDug/zK9CrmAaXzyFw7iSy4Vgx4y2kKLpTg+m0q0
5wFmV3FKtLjAhsMOZ/lN0+4QMoFBKKWJsWYV/yTWBvBB78LG9uvW195EUGrn
lG+SY3Zx5EhMa9w9wkHvJR3RMddowU1xrJ/oCXrgcxjB4HhC6976BSbxexLp
en08wr0eilzfsELGZaryePC65C23hiosIinlHV8E7h4/ztSMygducRFH2VFS
seSi/fmS4bfvNVv8qZU4P22L3TG6xRPUO2gXh0j6FK7qaL+ozmPqJqEBTesH
77w24r/5C+5ugXT7sEwtacNcxoPk8iEA4sMLQ8jygqLcdjzcGmE+STy+pZyj
p4UcE5g/Lb5QkiCPpZ261FS5NYVDGHA4meKgkcZJ7Hvz9WhwLHDNscPOfeY1
mcupfgkgmDnHncNHNzKkgFdtrsFeUxC7K5AguVn9/2YgaVYE/MZbbD8lvsxf
fDLXjc0p+8yZWFdX5SRPd4N5e6VyBSWm9pOH8iwXl1H3FycVK0/SHFuAFiF4
3zXXsycX0sxKeTa7BkhgsOYtCvcoIrxNusYZ3DKxpLRU+rts/Sa1eo8D0yHz
Sjlh2AVUg3RVkyYVlB1vh0xlY9mcBT0b0jYGbzBgD+XeUTlsANlrENG8oVgy
JnmyAQEtbjwf/ggYZ9Fs6j3Wvd56y3F3GU3XB2hfegIZvmLL2S68bpmjl59t
Zg32hsRpR1g4RlURVKgI6MFAl3gu89AjJ2qrlPAJw9vueuQ3KRl6+V02iAb4
XLO7/0htv2QLbLyhkVvUlNVPq8UN0XG91dpQEbTBWpcFEi7vyBIiGL+w+7JO
shsBoNWV4W+cpsqFoT5pzMxuPhG39WgWsCWpbiDVMZHbf02j4vbPUThFukdF
1UgNmwTuKHvN9dZg50xxGp4k+LhC5U3rxtgtMtxfMFqotcDQbjCCBpyavBCr
v2VZqew0JCk4+sOZfHqSZNILfrEC/pvWnCx0WW1huEgoby+H3xNd9zuVfG6u
ioeQaawnah/MdAzl1IL+IXZoTzMHCMf0AqKHgr5kRDlbNK00wciJ1lgSeNT+
e7oJhpdOaED1PPphoyoD1TQJa/0KCGo91iQOlQnsEYLaqKOFMAcr+vHmHh6T
DWXMiSnBWyYMivVAtCBkq9dzLxnaq56QB1GDahZfx4wOQPxIgZFbMwiy/zyl
VzJbNIR4bnfbTYn9ah+5T/rejYJjGGoGcnwxSk7taCPcCj33zpZ+ObOdDErD
uLFGhZliPqgnryk6KcXgUUxK4hoI9X7JnGlzx/PLRWaDXLxMY89qYyqkAgU5
x7ruyuvLLBai3tUcdOLINQ0i0oNgUwCQWJ7gNa2MurdwRXVVZtUDbB0P1hUV
EHuovHV8k7xvqdSp1g3zeXJ6rDV24yYUelClFJ4ivI1gT//j+KqUd0QrL2iS
kDYGJZnAhdJLJSiFK5Vk9o9sZR7mm+dej+d/GhPR1nI8KW0Bg7M63f9xgfdG
O3eZoR0UUBgg80l5b9pw5z65D2vqt2yJ02UDcBuRg9Qmqvzt8xcufQyjKLJj
uKyoCK8uqeXPg33RO9TuNn9vga4i1AwAc5kjAlUptUu4zRAkugwRwEj3BPt4
xMFYQQHQUN1NYlJzjw4zWtTp9QNdv+AeYjMOjdakdg5IiJIAYbKtPxIJZcYF
/3MnPlYLc5vfSUMFfvXYb6hMEOtCJC4VNVAiGM/LCzgkyHGuBak0Jii2AS6M
XSebUoCbv39nVaAaLc/Ytg405F5H6jTqUaaCabSHnLwj3qAMv8Lhtup7saXA
Dau6p7q78KvADo1QiE/R8V+O6xwEkdbDQK30ZVFQHU2HzhF5Brg69eDsXPy1
7TMZOHU3FblMg/5fks/bGpbL8jwJ4nMSS2u0etQ34Vsdf9Hflv2pcwrFCV1A
vVTH2nIgmJzVTYp0hqLSV4pb5kfFqbb8F3BZCzJrkasmCyHMwAYeENCEOd2U
JidGl/5oWAZ+YCOQAwxca0gTyG4iUH6FW0vk4m8G20rReli4gsDjBLr6N1FT
LqRNvvFPBUil/rZvo0C9yx+7wLvBP1iknofvtcL818OVXEkM1gM2Z2A8Rtzv
myJ8IBGzV+nXCrHhK6oqMoGOOlIobyquSnwhphVJcfq7mwQE4w0htTcHmkpD
1t1YjrWA1XqIbvD0u5aZlkAZ02qTvtVvTxYewoBsrsGef8WKiZKYAYcuEbBz
sLW8JyTpSKfIrlorH+er+uAs9HmA8MRlwcDly52BWJBPeiOJjYVmiCDiSSY/
WqHC/D1M7HMKdrQkKHc278hXpU7bv8ajHkBIuwtWAT/BFl9J3xVm3/ziMsC9
X/TLckAmyixLl7tF1/I6winblorrojBMpco3JSE5V3/dYwqmpftYvbnN1cL5
+vT4lSmg8wkoDc/ko57xoOn9nqPEzJxyEXIEkqnji9zgcnvxU8+WC+7uDP9/
gtz4nTqkTCKUXnVJMd6tnek6ZKypUd35DgvHUQXwDj3S5AMqJAjY7bg9FUgs
BceVkkjpEsspGyhU07kKf6j5maEzOH5EI7fbA65DRX09lRtjm/cVj6fUE/n+
enkumCXuU6xYj84c3zZFg8V0Fj/Y559pNmpyqudj+CN/kynarumtmRwEro7y
lIEiTDljMhcVV0sn5ixq9fDoAi1AzCKjC/qdGVhdjhydefT2l4imnyJuUK/y
9EYG78hQCo6WJ7QCOhJ0x0PEjm0cE4CpsiR0cjWmwJ87roLhRcSKF9WLyPuN
mHxmo9Qk9KuaslgVt05vjiUo1oFJkIhoO4ALBXW03b2yDF2NcVOJDCXqGEUp
ChagWEuPgcPmo++hFQ7zWjp+ABrM2bCN9TbqplKs9gxC7VH02XuOgkG65p1q
rtlDfeQ7OQEQHqdFIBLr5F0XVEogSY7JRGijaQQswxBAGmH7PJjewljbw3zt
PKBpH6EVGGJ5pCzkFhFxinUzGIXRc7H+9OigFjDX7XhIpcwXpl0NCxr+r7U4
+lNX7ONcOoVkjYADJsLpHqfPm8kr++3DKSfKKmbYm28GoA+mIQBc/jLPQygJ
F0hvgOrCdnBJwfr6WURehb/rHwGh7+9Tdi4+eSszkrTnvAKsrqxLZWXFAX7V
007ctavXjKaWvxrES7aaRnzUT24HL/XGOBGArw8eGByuCuAVLaTWRSNHjyjK
FmRWBv5oEREBldlS07hFhoxVskZoX162DO+244kB8Bdd3Dupg+u+McQymIIO
QCQISDft1bRFYFjR+FvLvzqQEiSt8yjA6gBTCzO/upWpUZ9w3WlSBePzM9hT
lQ3tvfFUs/PlGAt8gCgUcVZFFlim9eGk+P0XbdjYdb9Z8jykAMNK6Zx/TYqt
mKhl/iIW2BXbwa9sU4C/mL43JpGViSdPFMixcXOo3faacu+MjtisMMGLHMVd
A9AEi1bfxQNVvAuob9ZV88ZEiFX8KE+NJj32K1h58V+2XQaUXmJn9T0JUQYT
u9gOz44CkniXELyApEJdk805kTT5i1+t8c9bg2sJWfb2rfbaqioxcVEabUD4
Z4pO52UGA4MRpjNS7B4PUN6zsOOMXsi8bYENkAplwy1jY3eis6GQYPzrIYip
O5EFSkoG8dk/tVwgNnYHmSbutSNfFzFdiE6H4ef8V4YAb+KAcLR71dTbssyB
dWpl4lFTh+sBbmhqUEJWNghqS6ajsuerZ5zZLf5tcY9oLqM2QoGjMI9yHwSz
DTBeUQX7eSJ2Yw5cNzs5vYTgIxt7DuXSj3t1G7OJz0xew818unvVs3dD9yic
P+aa0FMmXVhcx7t+VeUiye5XMbV5oecp3lEVXlo+5wNQevkgP1wZ9i2KL4PJ
97DArymtwWtYhucBeyqhX/dqk3/yHljhLh212PTu4Q/XcHkbevVWol8aevBL
cP9YqCzoYcVAIotC1Ms7jv2pxK9gIXHMt+/TrjnabrRpfUK/Qn3kmkTJRkVV
erW+nIIewKoEu6+3zG1uMqAe8TKAqVaxuaPEHLjpqpoNXxmCWTHwtVMKUWiI
6Vjzev2TdvqV5XsBDl1toEJx7wbwtbUbvvfyn88LrGADxrVQq0wCT4fgLZ5c
n2DhyU+xK3eIGhknTV0i/pfWsFZB5Vjm0EINmfJ1g4xtSSmfAMpEz9DdUZYw
x2QHkq3427HEeURQaisEajwCwKPXaak5yFD0b099iN5gUDpYjWKHEU7VX1bZ
7KGgEL1EZ9cHipjF4ISxly11g/Jm/g2wfk4nYhuHDQ26+KvKkOBsNxLNcItd
zTg2EXhZC0O0YcW/juskin/b5fsHsft91l0Nu3RFQXqZJM+z5ae5NnUSi6pK
qqAJMKscrbDdqRkRLiZg8q9MDr4Z6ZY6FukSsGCDmrNjMMrKWGZMSTF9/abb
FgBTeI+VPf4SGm/2iYWqpe2JQ1PIvXPnQuhMeTl9yCyLqpfyuBUUc3gBde4y
MbEaoVArujcBUG2rvR8B+a5TUWQSlltTjOegB6TbqMoteg1U+bNCjOYlym8d
qRTzrJtAmRlMHQ82MGl1Sflk02kf4Z1oje7iSXSKMmMD91SsfBmEyjP9bGhv
nAvDkvf5K1BqtgVqmQpHf8VnLwNUxsxp2VKon2xxTzxZFgCn6AWyDv5ngXeS
MyBr96pYrQreGX969Mq+UeAmWcASbilhAutawohaW9ZjVkZFeJlr6JADdnVS
dwiU8bIi1TxwqU7NcgDn2eFm4ReTf0i1jyUm+NGp+XxXKPvmdZzNfaOeUHVY
mUMQrv/o3m96j99R8WtkHiOiiaWUt+jh71wMlqweskDvyMay8RzwzpOpJm3a
Xwh0swYHeNXuSLJ5mSmLvbIJ4D377eyfrOpNvnv+/cUulY8WmyZtiHi9ODPs
3HI/rmZ8StJFYF8kcupZ9Fzb9F9oBTLW+P6HX4V+7YTmKhMKSgRWG66e8BcN
z+1orbq/gxTjgmuJF8GdRRWtTfEnUY+i1JJzSDoObl+pgkGr4aE99LMlNrIr
mz+iqwHzt3XOLITlFxdN3YjEtR02z4w+tLD4SHOJZJcVK/4ZDTzGLWzZp8/V
/OOlS76mHuxBRVkA+xsHw9/ESOaycwgF9XrqeooAyvinOpezlbCGDjBUApUf
hMdYefRKYJIJgKRYcTHTIDsM1/qf9AFZob42ylhN9Hf13/MygBQRoROU5JWz
RZX0XFoPq60B5hzVlFP9b4POPfxXDmUqFwCPmPwF0aAj7B5M2ViYU3nokw6o
e7MyFZseWtgCqoAmnH4Q1J06xefoSqMSV2dBNGQhWAXfNcYosl1yFw8zoRQl
ozOidBHYveqnWHsIQTP83/FF5yn6QAyORSwcEiOtt8yJJKAu1ET4E0KvPh5F
CIvJ1QH2Eat3QIJnoBGbFX6b7kvgg4yBdtzBD8+yWD76DCMxSj1YHipl50Ar
2g8sHP2HwhHy8j8Ir7ePB28Cg9xQiZ9cAJD/Z3E2Tjmflo3WDMjpHU+Uzwql
T0zeRGLzBKfhdyZaiAw4hMf9Wc0jefBzWmmHN9w9F5SMdMWuFALvouun6a0A
dGTtVLpP5FvLNEwaPk+O9R3j033tlZ+hV3gN81Ne3LgXydeXdPsmQkA4Ocjb
g3wF/Y7piLA/eX1Iy8uRPbZv1QDmASE6FussAjT2K1oyLpAgtKFtZtfESxJr
DVmghHBBQk82157j7n1YkH328HglPPmaWMw0sAR6c52aDzd2T6tHxcNz4nfc
9QyRneSp5EDCP5gKsH+zKSP10/ib1WcAnqCQlPZXSX74WUJI+7DMTB78q6t/
Rb0ArCmZKC0mUTic+U1b6uMqN5jez4D0YJ20m1DBaDlXVjSeuMAHDrDpy5i9
b1QjhZD0Ar6e0+5d+nUqHKvW+risdznQ4XP4ldgcjp4ktGdnYwfZtx34XjXi
7fCLDgLVNuaDQ+C7NGy9tvbGdzU/crd+W8x8oaWpRjdzx8X6jwEetQHjTINS
/2D3rXFeM/2V4nxlagnduyx5wo+DrnFUmEKmaHyLbIgwfWvpGna1lOMu5JLU
BWeyWctrKBy90fSOmrO9OgQ/ttaTSqVkoD2yRtXsOQS3ArowYBuFkyJEswLj
kmRJ+3OSQ5Ff5f3DEr+b/pX3y5wllesZpCEHyb2YHEj3gyA7kPGeDgJBksQJ
1pFs+APt/SfDV6hUmqBRjpUvUrybVEYGLs9eAoUAeV5mKdPFKrNMBTkoDOKy
2jSBtcdsoj2prq4h54nEsMyg1+aXlDIr1vxzdDNtHBvzGV+yCb9SfRexbaOz
bputnDmsi3krnquIeYWjxoYdyuWtuxRqGGdEk5NDV+Fz78dJvFPuiCUq5frE
GK3fDJgPOq+N9Rdtr5IsvysMzy5gP3Jbgj0hXYQyV6agFHcMV4rTzbiZWSHf
hcc2ep+REM1To34NMc3Pn7mF2kFKzt3KyYenWda3HNs5QlzIZOCoMPwFhPry
PB/5IUKVTK5NHih63WEjiT7FtPXTUiDpPUwMHzsvclY5rw7jNSdjXCxRLt9Q
bLs+/fe3Gjjspzvuw1jTKcoWwDLhCGMLjAHzoWf9t9PuAlPsv+ogENh8ZArs
xw+8uE5WO6LHjzVx3ea6VIGxCJ+NohActa9f2mIvuK/wzc70mo+39L8d7KAf
W71bsgMdGYzoiQEy3Ar0DtZUk1xZHh7nHFbJzlu4L/ztVTT/w18Wc3PA4XiE
8e/EyVXJV/mKNJd+y7nb73IhzoySbT1i31x8YrFUcelV0OkgYv66nyhq7UTZ
TaFN9YRXExUNX7L7ZudbG/bHQsktSVm5ESTpBddWcOAWKaSVtnoi0aAE/UgX
cHHnf7eTQtZG1oWu+1Ep1Q+xSVPEv4HSA5VvK2GCeKP0uzAO2FPDxZ69941d
NBE9MLv4IIYJOf49d0eO52eo+MKGQINYMQLPaF9GFULZOvSB602YCAH9MtoV
yWcaPByk7ND9F4dwURzHXPkohIFzTKefJfSsbKb+/D9SRtUJtKzpIIJV6jk5
EdGNNZruOwyk/1b023Nce7w+EkxBaGtF4vHtQkCf+Fr8SO8kVQxnnutr6l/c
rhef3WKKiAyMdnILWsVIpLMFKwR5/jJe/KIShonFbD2kpA7kGmdgs8gZR5vO
0b0eoQkqq+tP94fGyDLEjgbLuc8/fLsgGJ9DcEGZyCTMmY2K8eTATh2MYj+Y
JZ/zQVGWoN/ln+J1cGTmpLlNBXdA1gonIL4eUEfPVV6YNFOznR9nIcPY3tz3
vECF2t1+VA3tBidCUbywtBp45amgZxbo5bmQe4be+CU7lLwv6wtWXDgTULyC
0lcWpL8Up7Vhxfd3qF6G3cE9t+ndd8T/014DAOIXHz7jrNYvbdbMuf01Vfrm
mmiRCnjK4nI5KVV6uXy1UNkjnJeXRTApjwMdQ3Si2GmFNArLAZZfbWylVeBr
W9aSdiuFcopJQXLR/EnLcZA+Hkzbu4IEp5880eCF8BgAkNGq0XpSEQuQf7I7
ez9TCwa1H/QAa8UDoJH+R5bv/rCeDEDZHJIS/OjlsdesZwTBiEJI4O2uBMZc
YjXYIPVODkVf5qH/zHeqQBp6fqUnddVn9ExlnEy5UyfdOwsu8SNZkBb2/j/W
/ihymmoDASiGmkmIhNCRx2/tHLEwAGar8kkjqd9Pn0i7WRbjqDC6Zn5JEIm9
VJWFMrr2jIzv2w5hcMgACFKmlxD0IGXgRU3aNjTcsfST1JUG+eBo4MxfXwXi
owxYjndWTOcHQsclMicYtkKGYDxvjqrxnUc+GN5F570PWBIsl0kRmzIaExDj
n+bRWT/d9ZRqaWpRotTJvG4sVkjMNx1oKHRu9R66pgRefKTKMq5vInCp/oip
O6HQAKnHL8RkbmzB7W9llk5uRgac2ES9tNbw77xkyt+eGJ7WEqQH3CtOaZbY
+Z8ZvDRCSf6GJtOayVzC7zKeRa2mlLX++7k9AdtUhoHQzZZLJKl23lvPG80v
rcNxt1ZC2YfXskcarGBKeC1SDkzN61x2fwhvzZYEA53onAAV0/DwsMZyBRT1
rX4EbacPTZ3Kab1X4oCo8+3jGO4YsNRRhvuwV1pLtXdojZh4Wj93kNejtPF2
kKLkfgwO3eqVgg8b3gXAY6J788o8cIrdiOl0RG69EZuMuLzYOOQSPycYwpVy
LuBVHb1yVcJkhHiRDxiZUcs3u9JpdXhJ6gvb6uEY0cHfabpCpdszjZ8aAKxk
Mc97+JyqnRk1waU9Hve7EsOY9sxVG0t7z0DKzoRrcC6FXs7jTqCCr0v8zlaT
vT7MaihBnJmLct/Uni+tkpHITUmlt5umNGzMRIdTXIVWoTLot92+hcMULzU3
WJA1WJwKg1wUlHF5KlCniXBXhazwzQDqn2BjTsPqCfUOBSJeec8ZpX5eODGh
XrvGRHbFCXsrXDzQE9TL4WFRpJuh4cF3MBsp5nl4ch3q71K+zn0FhAzMd+9n
YEsVUhiSJJphD2OP6zvqNVZ1U1nvUbV7/hvanslOlfxpT30sr62xGyfF8OeP
GpjT0SUGHd8HCNo65lzTq4ODLbjq6pApkdLxZyiv7wKiIlE7mwSjronBa4mj
xxsl5KiCN7frvV2ahVQn37qquR6A9SE=

`pragma protect end_protected

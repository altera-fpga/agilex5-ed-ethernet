//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VpX4+ryqKV58Z40uD/MUQ4RRAY/gTRYauUAGz5bUz2Ogr2jmZ7n8Ir2ZGYZO
zjGW0bsPGUY0kV2a3bdPVRlTwwPizUtV9ezuED9FUAVnEPCluUDR6TeaSqZz
5wpyeBVxEvmyixWNvl/N4a8rLwWrYU4Z5l1nYzpbpONTTWtIBL62F6YUd5V/
pmYH7Srx7l6R8qeT5j6uTXrpAxwCwQeHhDYDb8RD5Yc8Ua62Zktb9CLa8Qy/
SI26SqQ5hZU4k5BnzEiZRPEZeFCGU6IPiGhjb4tgmsQLmXF9FPU5jtu6Z3nX
2UgiNy+gPLFOIeXDohTVNNgHlMjCa7s3+bUYGqBZRQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cKDC9u5GEdxEEpHFh8S7wel5keGSMmurWp396unOPYmkWgMOdoE0cxMTT16e
ccOrKXv9wRK7p1azSM4k2TfVbMQgXTMAn5uX6j+Y3kz8Z7siXl7ubGIcXT+r
4OMaZYRRUfkf/BmJeoAa4oVvug9a0RtCbXLbe4S5b3ug5GOSiiC0KKBz1Ntj
XUbJGJfiwV8edvIrZxFVHYQEh0fjlNvMqidcD8W9mjVWC2Ra6e+35GVd7FQp
mrnUy6HIRwsdAxBFhO+cgF5552Wp1UZIajlEFlo9tCgBR3TT8bf14qFr/mW4
TzhTBeJ/ucuCFaAqpMbZxAS3h2c1s+atGu/vFOVFsw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XEID0kflTrGUv2tG6VXQECi+a1rBTq9SKiKyrTEvD181XQfyK/Cjkd+tBXgN
6tJKaiCqiJl7tGgGtyR9Q0Ihw1WhQNjkyNVDlOedMQ6UZw/9N8LM90knt22/
ZRgg1B9FCCeRv3KQIxRygjZA3ZJ61SBDkbQKXQ/C7YIR16UrnpBMyYqzhqUl
yQKwEVMF0yzh1wVo9ZQpLtqCvlO8aKhwBSblkJAvaiR+z20O7D41cuH6DTgO
zMskar8gQkPNmrAwgr0VaKgSW6K3iuUFp95czk6Lxip9i+iW4GyONWKiWhS0
5agZC0etnQvBRJjQZ5+iS9LKCIUEPaWubvEJbmdMRw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hfckc8V5B9Os+YaY7F+7OkFgY2Ogw8mYDoyTOyacnh6AsDg15sriSchov9nE
qAYRbJr/q0SGV20ofIdYijmc9FJmHqYPtMkYc7KzAHA4ecf4fnpedNrwVlB7
8i4KojGBRaLMaNxjt0wB5qd43q9QYUvtESaeo5srkS5m0kAlz7MT1O7McnXO
eiW8TtHtUVAAfppAbz76UM0SYXWOO4+BdOIA/6yUyGB+0UQOek0wAl52xU4V
3jvaHuvn5vXjwA6ab2443LFBp07feKTTHDYnE9e3xjSM/eLVLyIFolithWfw
/GNXDQAAxsRwAdqKKXVm7BoVvD1/gfUQ2cM7M9WG7Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bRY+pVZ/yEGd33yYCrczpLaiD4l9qwO85J9Nh8BdvV5KtkwQXbsTDXH0EjAW
PI8W/RIiKdoRI58cHv7kSr4ouVkKUXYsWjecSQcMf+4hZr8eKJTJCWxEKpPr
fGOfN2w4IRaAM1A2aM0r2o+Zq0hyvwfqyI/HsJQGXio5fPOWSJM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
q/+jebGWzGEzlgcLxGUpceL8fqeljosBOmWjbw3YTB4I50jM/psGHWozt6Rz
OLUnGHHDUc+yUqEFQMya7wU75BUoUeNLb77OY0YtAje19qZj0lnlo61l9LX9
SQhSKBcxTxKcqnoHZwhwyHMM6qYW2/gQ5yEK4WtNk6vgIq9XOKaIXaFK5Sz1
Rh3O+yTPuEX49/w8fjsBjvcEWpH3ecZTNbZqQ+DLcUiD1eTJWmppK5bpw+lY
7zZDh2TA4LjuFui7ti9fGfhH7kJTrYcDTFe50uyA2f/Vj+iUeM9XYoPM9tQN
PjA4h7SdJE1nhWyOA6thAKrLJJs5qb3VJKrfyRi5ttC+3ERydM30CJDGyQDo
CeYbwv2FvDsoc+P+1Z/OGQAd/+qYkclGGBfb0IrRtDDY5AoKEEhnwRdWXKvy
D44t7WzD80q6cBVXfd8fkYirKOXGXZR/0zhjgrWkgIicbUmCkQ7zMOmA7iUr
CiCfDnxEdDwkMYPbbLF5oY95R2dUFxOL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z+foK4UdRAYgraO6iMTJExd1EGpn+GhL8qnGPOWhZs0dWfIuZauin2w3Jv6R
+fOct5divBFAwwoz1fyZVMk0NGuabG/BViVdv0R9BDBNk+G4bSxR20VBdwaY
V1FHXFZdEP57kmVFh/ar7s8xsyW0nK7MhmkLSY5Y8koCPo6ipks=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hKOdZGh0ZVzAYFfyHfJ1Ck50mJ8RnB3KAB0WdKXh2DkG9d1GS1BqTchMI5yo
dJClR8pF4/Ui7JmnLQpLe0qdex2Z6+2KAW5dr6hMqUZrDG/WarkLc6SGUlo4
j/phuD6aaJEWbryJAoJXblSzQxx3HX9O5uu+Zir1GUfgM2VN5ZQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23200)
`pragma protect data_block
oIOOYfitwEhg5sJVdJKmdsGbx1ScAxBshWR4xTjh4iSxMDDJEA0xRAi2r4qR
o7fjTDSJjRT4UJBKKcf0Mqz8Rui3LujhKhayEuJoLZl68CCUKnUM6oJuaBN0
KJ/LxpMj0i4zMXb/tWzsVCJ7DP/KDYWNFST2DzSZQRqWZIswBOHjZwTrr+k+
Xw8/cUL3OreVW0Q3DoGjO/9gN6gGLw2+LrxC1tz7n7MJV5BxfUZabSJheL0+
M1hOpOFH8iWMjDPXyryr7eU6HxnLweRsLqxtEwaJXy5FmuCwYC4d8mLmMsfj
h7K5bVYOeJBXH6wIkAIXBTfbyLyNsB9Dp5KBWu8pVviUzkjjfbpTv/bHcO8e
VDRjpuQSTlwbIQG3xZmWR6S0NWaNprFpq5K2xjj4H8M5FoWkb1C6GcNv6YkW
VTdL5rvPtjIfcz50D+gza0t5SUTRmBcrpTnPjcQfpELum++KonKg5pogrYEG
KXVsDpS6quH0KyO4IiEbApkaqrulq734t0w5haxi2V7Jp5nT6RtMJP3xduki
C9ALwpRiSJLh1sVRPep+aT+2NDjsYkGlBfhnfqrCQE3ZTsTpJzTv0CmYk8iz
2VmGC/Uj+wuvGZocQKMHh9nkQWecBlgqEEHqjgJpk43eR0WW9T5pDare6vQ0
6yfj6XVX6BDaACVBI26P0w6SzlsrCGHqRfer5RSRAdmz8pvvbl4vrCvY0e+u
/CDqwfgWk78rUaVIZCd9rOYoa/98Opkp2uQSPCO1rirxAdeDgWT93mdswxdx
/SWzFqAvQziMrKAcDjMqlUxsoptq1VXYhMeWn5e7X6b5fAGwv/nGu1A6UHvc
f5sE01qftBWJROqIPwTx2v+6w3Ous0NEW+sKf5QE6Mfj37SCF7DlUjEobdjB
HPeY2jhE0PNitafrXBpPvO9yPc6VXPNKefQvfyEBX7tZ/KnyFEmEcVaIIutC
uc7MVx6HwHWVM/+i5vwxtolnU82qHN15sHdpY07hVFmTXXrCW94LXb68jKur
dWgcK/hVaj+N7lgja+RshX3q/OhNWprgAQjCgzm3DPI8YNjd35WKd0bK6Nzp
XWhs524kNsYF8b3MU0rz4Y9DhvmaCxGvUfuJ5Hn0snpPqv7RXB/LtzEL43aP
yguhcCCFrbUND8zKlEcnFG6V+MF8GnY9BrNV5xU2EKTq6pE3Yd1kiIGyPtic
KZKdcX5fEXx9uJ8tfug0ktdbL6DHnknC32ce51oOShlrQ92OyqZ1MSjNxH1s
TnmyWB3x3H5wzGymnx1g/qFKYf/3K8++K0ADq5WgZROIRN6+85/hmw0NPsSk
Laz0oGxZbO82VQVjtxZdV2SPUxkNgNgQ2z2Cg9DbwXUYxj9NJXrPuiCU9Puf
+1kRzha5ri4fO8Uoe7kXkA+D5YelS9XvdVKJ/HxlM7FuvLFGb/ArcnpLYlpc
WX5aoRK9MVgasFPOpvQS8DmMpUGKxKp1yCUQW9SiZxeFeoHhkJM9lL4eKttV
ivdU5ZiwqdRdPGFcJHvTfn1icDDsF+XIFUvsu06OgeH26XlyojkCLGMvkqW3
s+K3Nyy2NopiI8QWuf7YdDTKvjJANMWFu7z8sFaVb7DU0YuV5fvAAkUk6J7e
GZN+bOx2kz9NlL8r208oklxsBR63hFV7cDgieY6XCsOlPuMsERV0W5g4wjcN
Dl1OlhYVz9WM0wXZ0KlHl3KTyuiurgzA9KguBodYvSqJu1R6cN3sex9GX6G6
ESPP6j7JckeBm+TvizayIVx05ZxFr0xjRPLYboGamtnUB5tMLTObmBbAOf8t
hvMJMCt0hUvhOCmkoEZb8wRmDtdIcpRHjAgVZ/tBANp3T40ZZP5B0b2VbUV0
vt7RKbMXXKzB76gDYQ4Yux8xdYqcWJNAogrYFreflBGSWMqB1TxgLYVMHPka
D94twjcx6r/wIaH18Z/11md+Lnz2M1DCoX3KGF+jEa4WhYtx4ZysRMOaCV4J
UKOEvM9XTc+1ITnNyOxyd8lC8YnRfWbirq0f+94zZSqZ74/tqp+vFmKf3iRZ
NV6gg17p38EkwcjdQf9A5S3PBEQ4R4gmlg/m192QT1iUBp34hQUFH3OACR2z
P2MihWFATn/Z+hV4KweeDNYU0yIYnoG5ojMYx4r0CdPnZMdKQWvPqAAzdjIQ
LHWeP+EiTv+D9+mnQrUyDvKwYhojePEuPqBXLUqAkxJJ2s37ES8o8ibd7cPs
m8dKuuBqdt70O5ETyibS3Jf5e/ZUzoJ3hPkO+R6khy3W+pJG71MvDhxRDe+B
UQQ3obOU92+2eZNslZzVOB//zjTyMNZDi9OtD9kQFhVKMd942lT2AIFg1/Xh
07h1RGnXiDOGjsDd28nECtzsh6n5ApCVYEPjliDx1gWHLvvUOKK64Y+DrLkX
/4423/VnSuS1A1V6uM6glB7MmsDBvQq6epGwI4Obkjco2PskYotee4Uga2h1
ccmD63DUSX7cGfrdAYu2eoQs/VllHaI+tz7t51betIFO0lvbfKkuz0TL1EQu
C4LbtIRGBrLgEV/EnWIr7KWWMSgnN+tnAt3lmwjSz5qBg37UCC9/54QXsUuE
QrD+TlqL3fBh0xdNJYM9j3PgJg/tnelganvEQjZO8kh1QV+LCoEAXrsySVsL
I4Q1TFNnF49sx9dV3dVMHwJdz21ub2m3d3u+wXr7UAOntW3/uTGwYR98mOEQ
d5UKZNOESzgoYCBQblVKMWxE3EkrpPCkEn3dhFO1lIapO1YzoQ4BWmjcAcnG
qdnsGVQQ1qDnmBbRwuQr5h4is88Km46Jay1nbArg0rA/3+K6kUK69Ff9exqZ
aWPGuchhij9+K92c+O49XY1ftGGlzQkjOsnRP/PeVoIn4kelq9SiXd4bLSwe
hGshCF1xYdcQ2GdL052HZjxp8zSfpetPobM4j8exZYJZPSERAaJVPtZY3vkA
R1Da84ZhVFA1UwUDqk58/THqIKiZ9SDzUowAwimGbSfFIwtekiTfokD6t+DL
cBoz3vkeEuPD0EF0IQHcMbXpnYNrW7c+oRnkdJBX+F0Z6qXkPvLa9QlVkx9A
jhnX/lNsMqtoAduUBLTn++iULyYtM24Xh1lOz1Vc1FsO/BQtIouXr7ZVlxyI
6ZPQLvFCRKLEbGavCAKcDurTZVWGjWaQ7MCcWs7hx7PiszPXWOOyrCvRXiiK
Gj89jr6y6fxOHcHrtN5Xl0x9CJLpMU4456jEBP838P0FkGc6tR7FZ6XWsk+r
gcpingrkuh7P/Sroj0nvn/FluJGJahSanbTLqKPungJ0E5/jNiGJuRDbTrKs
AdDbjaU2YD7TLJAOIwrKJGZ7hAbVcGUuMMpj0D3V1iLLDNijGErjp8/01yVO
NAE6MdIvmuUY9tiT5YzATqA6rQKceMwinagf8ZRBPm2fd7gV33gIcOAVsEaN
SccJZC0qVpL5eu8oBUZC23TaDZj/svZalBbOtz2XT/3TsXD5gIlRlC0Be8XV
t+QHk+H+kfa3VTxyJl8/2uWAO/s4JwPIcLCxaLJH+435j5Km/SLLu7yDqiCj
ui+KpqUBwChT7k62ZbB2znslbHn70zrNY9IEoYJGTkGkNBEL0FLD8p6fVtEv
egLssBJbSE1F23rFQQ9o3kyf4znBOD6kI+DRdcpfh1e1V63aHoIN4AAQxoym
eShA+dGUC5euLvygTGh6qReREVXUbKUgfZ8G6AN/30sj6CSgZn0xMjsu/YGd
WzHRdicT42Mo/vuSlhOhFHhh4KCwaURUZystmLlgEOC2iMkro4pOs3s3t3wc
fmLZI4pQmiFAAB5v01/3cYoXT/sJNvZtp4y4ySsP7jAli+3fRdpYvaCcQ/w7
E3vgQKp2WT96X/Zofuk7hcZ0a22TOeRmWEzUnnYy28JJ7KlvyO/1kgldxBgq
OCeJxtoaafT1QuOa2B3EdaEw1qGqZVIE2f5hfxHs5RSeJxA02qF6bWIGm5qu
wVMQz7YDHJ8Rb2cQ9DP0K2yNBhIdLHwBQc/QADS7zBLxRJe9g0AVPU1FMw15
mHkOS6wbKhpQ35QZcr87luclCRbojUuvYetHC+qIk5jKOA7oT4gflRha0GVH
EzOYTKcmnJf50OKsGBR1+cWsUBiE2x++7TEeztaSIxvaaO0cU/33ymY+XQzC
U2DIj4dxlRy7KFX7gIdotib7aKjH5vJ1Em5y9dxhIH0eHivt2wqoi1zPQRkl
CT6SxCzG7L4De4RLXR1L4ulo+NqrXj7ebRkEqJlPp4y0JDdBCbeUAJ18ZgxW
VqqlIJawcJ41U5bAkEUEpoR6MOiKrcwUvJpknOfaNaqrL5tr+SsfpgKCj+aR
l2RhPT8QDkMkTwLOHRfA/zxld854iwy5GIphILkUQ0b9ko0Aq52aNY5CorQh
dedisniUulzxVyqL9RuDNzv+ldXPbcWOVyCOvKm3hl3ArGKrgyHc3WAvqSZF
rOikvjvvAZc9m+W5/FmhHnNpqdrK46o6cnmE+3yPhlqXaV7Px+4H4TQ/Kup9
JxGrPHjtI8h+I5i3OMSTTftA7wgOq9wOCRBPYbSGS5RNkvPI/r7UmvjG0uXR
AGW3yG/GggR/m1qKBKi0UzspGc1zJAUnDUpGguaPKyZw0GkFLhv18EVb6bGt
ixweGI6b44VUVTlXLrwCmiCEHFxk7Ns60cYAwhLJbmOqKGl+WDi1VtpCEUE4
tLCAv+TLzXr/zszJof36UObJt2iw8zHSx+oO7SF8j6060V6YcFjoac8E3h55
sHX2gLTgiMZQ/2TLerMwtoCxI4sr/y+fOyUL9DKW28cIl5NaqMWNeBKlGVzW
dspbCckRkIV62tFNdXdKZGyuyQWyoSRvpR82YfZ7gYL0tq3NLCS1uRx+Y9hE
w/8KAH0C7WkJ6AwTELfiaXAhy6r431qVZUBcBQ/E3HZ5p3gIm7iIN0hnL1ol
ax0JT8zRYudK18yW769n/mVVVKcOZ57eKcKSZCuaERFnOYFEan56ybTVI1vr
TXcw6kHKRZGG1pM+KmnaxBDlO5J6dfX//g4wLcHcYWt0MOlg7kJiJ+jBLWTW
GW+jQDWbGrjb4aTrqVgTANsoWw//jSr59gAM5CbpRpxrC4aKZiSBdKw3a//i
i8DDsrTllH54uP+I9hdakFraeqmOP72fnfFH2vORAaYxpupzYjA7LT2iaUS+
8slazzcjMR/ajFfM6vv9Yh5BKo6HqENeQvb9bRA/JTZZiGkOPK89dZ2qPyuR
VKNgAjygwmv3tnjJ8/6u9BmTRQv6EFAfSFlfjgc5f69R4VLzzW9SD284H2UR
xagGB6inBkul2nHZHR7NQv+HEYKVL3+o2zQ4F2JZv6VTyd5eEu15rGk/oa2S
1YK8PF/Sbd6de5IfKxk/+AmwPcrCTc3wCFn8Bqva4s4IsasbY5BpnzA63Zcq
CbTcJ41Br6BcgAZvdEoovpsxx7WpUtN9FHvRyL5pcgaDBrbPuBCRolDp8n0N
ga+08iKYE96kILQP5vqdNds8YBnJtZEfPczCRA0LSlgPt+qe5eoVNEsXnw3K
I6ft8u+qdeMHGdO6XMttZZk0gcXAG3YCfBN2l2Fpbt+40n8YGik7TkW0ym7s
aJcs/D7RynLBssZ8Yi37EMztiMJYnqUjj1kQLJbfXBX5EJL6k+U1IPSvojc2
O03VkS5kkKo7SfmJIC3He0rfSPu4NQAqyDZIfz/xnqrN3FYUl2xpfeEQKhSM
hLNIPAa3ZrO9w2xRo5YUubtsLCzB35JyWOI7CVWZlYz9Mp3MkquUDQl2OIW4
uN9MNBtPskHzaMR7olZ3o7Y30GPD80Tu5TorhyHtvWXwawgHxjBxMU9KrzBv
N5kWY4zcqQ13p2UGj+/MdLjrzmYp+AggrSxKzc4KyR1AILQDlqQTxkW+31mS
k+7+ZztkhawGF9GlyNjkYRT/pd0HHb9wHY0dLu5EDJn0k8jK3gNro5bWYEbK
r64BL6F/PGJXq6tqM+LsvHB8K3zqvuHFACKSlmuo+SvsSOH0UwQLmaJRchqK
RFaqDDnpg0kwimGpwVoacvcKZVqttsmUE/nMiZ5yZbfWNPFU5ZSE8fi447Wu
SMiQL+kL5hrt9AKChg1Hpa3mE/CayUGqXTxd0sh/WNHo9AaiPz4n8pBwCR9S
//5zPDDzCr3QRCvyenPcxCDYWgKzrSTmKHhS3Unvwa62D4nYhNP99mmIpVP9
rDpWAkJyupbdERgPRtBITU8GKdpJvStfHBhT8IAPNfXy5+Ew2c2yKrTO9mlL
WeRGu+svKGRpI2uAf5NstJA0rP0eUYydA91ULFoQW+MNXfG97A+VFvdDqM3D
hbhcuLL2aN66dfCrLpkZsphwKVvBGesjZ0y9SQkf16qJiLIWTrT/dmQxbrFf
8+snOKcX6TztKWlNZd+mmkLmeji7vjFXUdEZtN/J5MbEtt1uB/TSFw1dfpgA
ujXGwjJIeWngNdC6gVTp9sNNY3ylNUBQIB4qm7LbzDGwOLJpL0S9qf8rDBBN
x9pLcreIDtSrl2e6UloANHnWyy5jGrKWC772F3mrLyCfEn98Guvd++ky1j07
BBKEwAjOl1Kj70v2QtM2MyROCDoxlESnl5Y8fZ5U54s4ZHhXTLNw751POz6Z
8WhN/dDBj+drtJBU6BSWimoePGq9YHldX9uJoNqkkQKwPFlKOf+Z7jIlVHej
E5RlzLsxw5kA3WKbdbB0m3aNuwzM/QJC0AECvEb4MAvZuL59zaquA+OqVJQ1
/PkhLVd7DLQsyVXxLZj5RUmVeC+stioaKTswfSgwjNZl5Zgu1vPkWTSTOcw5
33eaJDCTomXPc+pGHv9e4saTbpl4XS9KlT7Yen93W1cWzSqbkM5ATfHX+LFz
DCFG6wIuWO4e+Xrnw+knfdUK8cezvghRDuQL1HkEpkPg9a/YmPZYXQEDdb4z
jrJMxWeDqJBFCfiAERhbJi7pScOuaGJ2L8BZjKqf0y/N8JQTqIg1x0MsEW3k
/ItY+ARmiSFezGhtzGougu6dQnu/WhdxksDDPewEmKPxa78XDqYMe1BcrPWT
UK/ZdCWxqkpEdaTXpAQcFWVbnXk9qDEfewiGVepjASV6ATJjS0GJbI8vF29g
cUZ9bjSqdW50JaLp2AMH6Yj8JyzhgpgBhaPhjO2Sqnh4MwOcGF9CRwOx3XFr
y3QT4FjfDGTgFOgXEpZVBabdSz4PPv6jTwwmfviTD7WnjKzkFe6+qyfjHWFj
o1okOEtg5mufHkuwjdll8LDXgvXzlREIsmqR4UfPodBDLTx56xdk/MnrgWcL
RzrADkKoLp0QBiRssfMmKvqpi1bavqIG8scC99yD2aaYfH9IzqkzSmhckWp8
NVq7bkGQCijWWdfkE7uiYatjSMXCX4OwbhvUZMhU5kllDfqLSnMN6Rtt44nV
LnQNtqh0y+wTFIAKeTIWbkRIvfsLsMh+O2ILoG6g+7lsrYsgm+UwnrEnPPKF
aIm2I3huDcyEdH5y69xMG3z81z92BjodNrstOqhlLYOP8hkJ90jNJ0h5Cx2h
OZb6KOMlIXjy5D6MFpvEoRytzYskKOK2OCTFOSEa7ZdAtn/T9IYQo9Bqcf1x
e5B4Ky4qti1SCnB5OpElMPGRSLUnbEwToillTE8I7t5t39RRockheU/NktDe
8iXyEvsNS0EA6zizNH1em5jTe7Z41awJa8u+NQo5D/xfKg25Kvqi+BCWlexa
9Qhrh536twLZ7+TAMLewNMyig3uJfbqm6oBW4+k0xpGMxukMEjR9eHtUuDRb
HhAhBy5YBEMr1eYU3mMgGGOD3fthrlAKIv9gjCrLuWnTQ8u1Ry177QDMkhN8
gbTVFoKmwjzik0BWTytG/58iqH4NpGxh+KJQFIA+QDpe3Uh0YPkEmlvTkcJt
KCXJVH603GJAx7Xy6dS2YaDPx5UGUOgCuA/guaTUuiH/C6rCeYyo2Yrub/x0
j0POxkfv3xP5qLbI4WUeP+62ONAFa1fO+XMqgUBy6K83kbfuEFGtTSDntTjh
tvJT56ERc8vIdUs1JxvQGbBYTv4Sda0+U8ipzXrAjkOYwSvCgFAjKY84xLmJ
USBt1ZQ/JinaAPmSp9hZ1KYkW7hvfea+YuGTslYMjAtpPnzkkxWiWZsZ4+Mg
7CGxp7ouyAV2qBnPNwuhYtpEpdJFh8jueAFyC4IIuL9BP6XG0UT2lvc5lrqx
oY8zbJiDjY76sJP9fnpm4v3L0p5M3qsQ+uPOkvAOXO2V7o+YFpTvZ7wVSkZp
Ai3LrcZGTeSKddos5zaxh996K0C2Uu5LbiTVDeQy8KRWTv9mzhLLC+gY3pdE
Qyd57zsKMsRQBSTNJ4zAiXzRPTo/zgatrv7cuJtFTcJBlYARebVTuKP3+rDY
48CE3XHiO3Os2qG9cle3phmyIOvZWW4C2EoFtIGyuMhCnaF1kQBYbJZWG1s0
PXASHZdNN6jkLRlLj8Ui9IBi0FwiEDUSEVbuGDb+pzc4ITiNHV9qWuBRcDqG
xfCYEQXhNE2C/LtBGPuq3zMDQAhIMuD154TUQCfNfXQAbbY8ffmetZqTip9Y
fwxSOxG635eomK0ZBQ8wDDY6e8I/CZaZIHPVvW+WP/y8S+OmCuIqU4A+NWsc
z2ZdDI5OH3jDpoHJGWv1wGGL/VGcyDgdoGfsmXQC2LtZEuWTV2JfLsjBoh5R
L2784MK/LVkLIepjsDtfpRy4MQ3o/qa5Q8/rtWqRKhGWk3zIQZ2e2pdu9OR/
a+q1AyZXTXWCS14AKPneAPw7V8xqD0WM8jmP/8PyFBa00dMllfwizIF7eilz
5BdQqkQkbC7GfR3Y+IGGRrNBziVgvDgu6LDuAV0MxJluzINit7mSOtQsGxnL
t78jtkONr81AmH/W+b9voTGGAuPp2qdxrBcTHEXcLlFiC/7tqbKJzZYqq0fC
Dxjpn7EMtHNTk9wjin+CWxElqdOpw3fNrvLv0j4jjrr7NB6FMcUPN/wy44+S
Lc5fZ7Fa27GekG4Ke5DA5JW5UH45dBHxDHzUQCZVCZjh4hqf3c5P+t+Kjup1
R/V/794xJpy6lgAEVIDHqID8m/R7GIqI0Rf6Dg0EZnx7+cVMwLIhw5C95dJm
l6Y2vHKV9d5VUz9zjL8R94opUqmyvpfegv+sBdTDExtnOPj8VdbKxipnBpO8
V5FdaJdkRTrclnlL9AFmn4jCeNk3j+DcXt/h96RrAZYnXzFs+/LiPqwW9+pv
xb7t54rCSmA4SN4ttpma7RWinaaBLEberCuHRKR2JeB4y41VQ20dfs8o69F/
Jdwk5T539GlGJvYgPwashsbIqNDTEbX+uxZttliHC5xH21afcMpMQKI7ij7l
wdYo3Z2hA5mj5gYxzfipybZrm4vMffEA4rPp/wc2hRv3jwSddYRXF2adt76p
yc4HG/58sejXR1uMp9qTCefA5klB+dt/VeB7vmY3OXPtc9isPnkhi99t2v6e
8O75B1vUfval4iEZgOpg0FtJw3nJh4mpJBO9vjv/irmmtFcynDwVumLV6XIz
JiNF2z1Qrv9JGGrvmzwlYIoUMig/qWKXeRygvwWd+0qpfUo92/MQ30iOj5VI
o0rPK4h70wy8Q5rfK96T2evEaf2+Rq9scp6uF9OLUjp539YgcSz8xL0TpdZC
8yUB9w3OwbcIv4gV7jcn2/hEIbmTVrjhZZ06EEDp2DYTmKZS44FR1IS0jFLZ
fa2RHhMKC440p3uws2lj68mF5BntztradW8K1TILq0zJfMtPWIc5k/IOEqd2
xPm91Uzp6dM0EDG8et/hBaUAqSZw1xwxm2qKNxDnmgboL3z4tIffIE/HsWvF
VxwdZUkCqWmxUvXpjH2EhMq6iHXlxTws5iDgQAUN6mn4GM5/Dx2qdcKzHPtK
7PmTwdRnIuH8snaWO/zVt/SQDdenEiki++ugAIdDmSqetADrKYE1C8N/y4jb
sAj2spAbxJdcpGCVZOs+ekxxRDJqpY4BRkCm22dzEdXLXeuR7nGp9t2tlOhj
v0youvZLcEE0026SrrA+POpf0DYtXvuB4NsPJ994IELtCYJwHshVW5IUd7eQ
26eRRJfz6YBi9g7jrx/v2GbFoRxlGUn1y3qEPYzSc1c5D3lPX0MlRw04i6lj
8BH10PG0UzOLe6PTn2olLYrnD+jPQLgWAL0DdPUOC54OqdqNPPzJK0dyLY9F
YJ60QdbiAkMlh2MRwi0zVlDdUElAhvUN2KlNVxWy/neKW+FOEuomJEFdksmv
YWdnQGAPH2eYTIZYA7IS2gAgKblEwuUROwepMTDmuLZDDtrsxXpRXKEYtXyC
vdZHkeh1NYNQwuE/sNqSCcWOHe/Y57xCEc2ITt0xznvlhuLoi2hkYXzGkYaP
CYYAySHPGKeIDaVcssGPYD1f4Jj1vxuBB3bVcAT8PU72DMC++1TQVGRwNg/4
n1xV3vAbift707g5eMhlfQCsZwXlZA6o/U1+3S2WxFrtidFEg+60SEhEkHfN
qtickgpJzSj5nKPJ/WkR/lGuTZI17HyMRMaysxd7Q38eeK2mGVwB7UhTJmBI
s9gG2Kv6bsHOvYxZiwKGPlhni+2P0FSnpoc4/6KsEzEpC7j1OMscJCnvHNJY
RQtKQ0jFdHu6WgHFh0nQk74DdNYqMhhhmPN2u+nyaOddyZXwIkSlGM7QqHwI
EW9BtrcN1BBiX4eKYulzUEcZGBYTN7KfhcHKQPFR1Mkh4991W+kIfZ/jncj/
vre19GzPZMX1ieI6Qh1dn87p5W9eI6jlxaVwj7SfXZKzpPrS/1TvpzgxFKL5
EpEodfmiEBC0z9rqTJT4hib+glxCacpu5aKZpZYfD+9Vt/IkENwu25xLqOz1
340q8DeAZc0nQrp1xFmjOlUDFbxkJJzvSi9Xj9M1p96jZHgugp0IY+6mOSpL
w3qIJhrYuZogyJK0Bnul5O+yadtKAIfje6mKNN9q5owLPg+hF02K3MGKguUH
UhiflkwIFIGpGdyWueu7jnsJrNr37KTk9HFtca8fTjLvYQzYGULxfydrWWJK
YpJUx9d4iQY35sPHcjjWLyrUMBqwr79p4xJ4seztBWI7Ritzb1ql4Okz2PCy
gv98n6EdcdnlwodR0epGJlQ31UYQL7cy7kLTUH/gGRBR4qC//9g/00XwGcu/
pSQjwcOEbuI8ipsZVWjRYl95KQ+i11I+dKIla1bww4GXc9l3z+6AxCXkdYdt
Q/YjlmYMoFX0f8Nu2zR1ycXIuIswbbTMcjxmD0oLJG5GZcJi+UoEbiyPr/f7
nFJN9crrRDO5qetNA7ni9noHXyAe0hLgPThYLUmhGd4cFVabPbDJMLc2cULG
UEx2jvjSj7BI1tK5w5dCMdrGW67aFy9PdfsXhqU71gbZXH8fqLLVx0W5dBo6
2xVMFe3+sDRrfvmA4DM7D8R6nX+o6VaD2XpxEvS++Cu/XqzpqY7ULsJRSXQl
xGD5qUPHTMEvAZU9hFExw962WdYnRDZhagJbWWyV6tscAOvR7sIPF/WB7ArR
mXYz4DBXo8uSC8ZGiB7NkdW8/oOPo19AaLbGLBEjtbwSdcoBD1UUqde32g2K
Bnla6lNQFYMxTyP9ip2SDhpHsvzfRLq0WxG8ek2Qr9WkOhAa4n6rKIaGCHsQ
Ho/c64wSzVAMbcLnHk5o+UGkEtQrxy4Yu70zyUiXMtZina+eZevwM7ckoYFu
6K1mYz7HHgJdVv0630OyW+TRXTT7C7PV2V8qfPqOcdBLYqX0pbRW3Y6EbyUf
pPwPhuQQE/DHAV4Qte9Tm8RWgXZdZj7KBnFDBdvBNPPlpi0ZLLdKbXNtlqQQ
kX/XTIDxbSKanBvkLiPb4aZaF+JG58Vu8DodN1c/ySgTRV4pqlcis16tOoTh
8jzXc7UA+wrrBhP95Jfidc5Vn4Qg6hbPxMAFtZUt72wlymQGOZavJ979b3Fr
3e2t+UJaRHwZlnWfzaA7NkW2BzxvOENV8z0n9VszB3ySvO+/XzaH+8WHfzWL
nrW5R+mgwSnp7Du0Fpya06YlywhmnyQOw/lNORk3OfrocVUziMVJUOFv48ls
1iAuAHGFPHlam+SKwkYD6A3DRezFfY1Cc9/ePb9pwJKEtDFarUC7CHFXtkla
YEEL8hRo7LSKXLJSXMmTJnJYZsx0BSAaT1EJCqvro3M3igWMIY4nP+s4EzmM
LxW6Y5Hwu58sXlV7lNGo9LgUqggD1NtkLwfvOejuyJ6pDhpuzysF5u9IbngJ
YNHBPvjYXa3zxtFT1mAzUtjQ4H69/bQYc5ScnGE68bKzNIqlSkjHyvQUW/AL
y3jWaMySbD+Ga79agZFSm4X4D7zvDbx7uXAdDw4h0xZrx4mEItqIuualaZ1J
tYKYOz7gkPX6j3+Ql5qVnp+ZpAvXPne7uJdYJm/JGZ4FK+JQ71D8d8+gKsWv
F8+HKcneFrxO4Yh45KnGncuDZZlJj1WQWgBlO3zb65IiDSnv2xW3hiTa6ACk
FJLSJA/6QGCy6PcPwbUp29/HWl1y+H9br28hA5907N1S2M5wzgQpOXxbkWnc
ArCz7dI5nLlIULyZaj7qmWZzgDvR5NDTv58xXpEqdCkiZERIDsC3LcAf7X+O
HuWVDqt/KoneNxtxUbpbRWXuSDLgjquMLQzWLySJ7ePFva2QXT2Ltj7rlPCR
3IqesyPTSHGo2oI2ccIgR4RhmTDek3cTP7PYULEt7TER38brKWf/N1il/BPs
EyVq8RoNg6X9MseVbuUl+njBlk6PROZkAcho1tSWeuajHh+yVOiIvhSGn1M+
Db54lmwVU8ZyjujvKIBQdP1GTxteWP4kO4/PQhsifTUrl5D2CSMDO1w7xmgD
2vTiU/tORlVsL3jQv49FF/Ryz1/3XYHNknyLpK7pCapFixtHzkiX1oVQIJtG
7LjGfrrHZ6fVNeJUSk01ZHs7n484moZaqgrYJURDQGp2Gdf7SGZHZUxaRnWz
naicvE5hEVAxiqSUb9LDw0sGzA6msYWE+dqoyW4nddVTYIj58nG42+cHkt8x
anU12d8DConLUm5MglBZZt+aq0k63YwNyGDFBwRBKe6049aVatopLA6ciZ5b
Q8A/iaiBfTT1P7/guecSIKZYd3uLxY8SD5bT40FVHYfjRRIKv3Mu5b1dJDYD
YDsmp0AvGgkp8EMhmJ99vxv8YFsBfLTtxKKo6Gw42V2kInhmgvS+VGTILsu5
Mxsrd4QVeTnLocISO2RT3Olih+bDqifoLuXZI0zIYjZwvSXoDAlAHm7fa8iq
4HdYKxibYqO5jiCc3+K9NT5PfTkMioHbqHinHQ9MRgY32Yc1w8md4ORubENt
CdZm+U0xCaSdu+hBidLXwy/gRIvh/YSKDz8cuJ9NKyPxt6bsxUVDGMc/dwlQ
SQl/AaVuN2hM5Isyj0yt9bWB9Yez6KJHaOaWY03kyECk580GRHAK36NAEF3w
Vv53c+8aXOY64+l+Ma/I/6GkP6LeY8s24/pUDNJkpFgGm1ryTo1Vld78lkZf
Q7AhpH+PqMhgK3jjJKhEwRACKr9SnEOxxRpa2dJXSanOwXJwDSPDYQNIR4T2
MppMXay4QWPabC0RP5wBn5C7gKYW9heJQBkrIxtQE+oWFDcJt+u4u20f7h59
NjgmSPtiWq5IWrD+c3THvilHFRSWibF4v3ksyJzGPceOGy//eM6hj4hZXWPI
bDzkxQtwMgHa6Hd0lvOjTRjEKYmsOTbSlb2WN3mUYBEfDEmgj113hP+0wjcs
dsqKcdi1+/MFo3N6SM9kBJ+rK6u7ot2Aj5h3Q1GcoXWmzyZXh/Qw6klrZpaE
7DsIOc+vpvbrE9MPEu5p3K4X57tWbKoWqEV6WHbMc+zeARV9KrGdEKXwaC+1
an8RCUAN1LdPYqa+hKEh9bxr4RDU7a/8B4AH9GOdPSwQRBwD8nuL9QPogPzJ
ktCt0bj+cPL0sBbdBCs04pzqaYtnzeVWw4tR9Y4Jtpsy4vdg2/Zr47TfSb76
cTGIZepEAJufkYjRsWmqMoZYjU0x3BCpvNV5xo9fF/OqA7csBLj/J5PJSwrc
qArS4YoYOfh8hMDGXGRgzi6CbDals38+1lDR44co+pqrlHrhP6LnFcQWxH/4
FUuPZJDJCDbdBu4UkEOCL6nDA4C3GImSfRa8oxg808hpf0dSiNlfC10IQWge
OQzQdVysup3AArWyRqOnpo7ITLJuC1iCsy/lTf8jwtZKL2i6h4GAlSf1gQTD
hMi4lHqszsnZDbNpg42a5O1cKWfd2JpkbbZPQ7DOGD7W3SSTBcd4ScVP1vJE
jVHNAKsi80Us+UGzSAklKX2lw6IfOfJVepjvvNjG0XcgXu0oJ+x7OrrRwQrq
f1I7fFn3Dods5OgRiKE8exeFfK9hZNIt6dpigDkbX9NNy3tkgPUYu5ygBwEU
NhDjGfuD+5q+Q1I6+hZ4CXa3qjbTcVKfpuxHNXR0mJ8rqibT0i7/vGAepPF+
Md8+SpPu63NNvJBRIVj3Xaqs1Z8m169NdRi5Xf/woZHmvFlcPMkhMXtjtnOL
myMYOkhRMkCok1VSGLXl1I2nl3H7aHqe1a/vTGroPJfSjebfcLCk04oR+JOU
4heDl5gorU+HQTw2L5i1nDgoqDDpSq+Jyy1fl73KO1/UEMxy/4Zj+lCf5XDh
f0MSPRQV4nFLymXbhKjVpxSbxMtSmdAaUDgm7biTpeL8XEUKVEv4hcZaNZB2
mcVNzZj57Q4CzDVExVMKxCYlijwUiZpztOA92GpQ6GTCHL72DJ/WiziyBNKp
vA7ran7+1gXIxOIlBmhkBXPndscGSTakZ5cNlRbFgzD/NIE0nx6wGSVB7oOl
VZ2cRcXk6aTH1Eh4UorH9op3E1iqj9va4rBMUSt//BUKIc6Lm+2PVn18cTJI
0o56Ha6Rm331t94NZQxhJI49WnuH5SX4OMqjBMq9YNbNgdpoA8OqcqwYB8wo
cedyokdAeZ9k68RXSrDn3iQH3CqmraK8iXPPogD8R5oY5kspFmwh5jGU+Kaa
olEAp9DegXiqd9MvZR3YYpbyDUkgbCMxmHCzsdNjgJU/aMR46EldOMIindQ7
SG724y51FgAKZd3rLRe7wkU8j7jyiGEHcZU37Nv1UGBHFK2RoX2f1C8RL5VS
PMqiNhZwHRLDvb0AoLghhrFU5J9eNSZPnUGqovV6/7HVi+gaHwPXTP1Cpt6U
tMYCwVO0LcWwxpmijWDH0vTg+omPDKzPQ2lINCPFAVTJNlChV4YH/dmriReZ
HQ59rb/yPfxVOxEVSaPHduvUi7/LcvYoX+o4Ti9xZJiN+3bu4hchTrus4DIJ
EAkPV8J+y0ZCy5LskwdzugvPUejfp4RXmPvQ+8JWl+9g8EZUo8W5ujY2vz+F
TQMQ2GtEzLbK8JlkPN4X3HpYrvRSMJMJB9lTYQJ+vH6EjbMedyrOUXHIZG/+
6v9IHB+l/Xd4LIJHUfaiXliBzUZQ//h08rzaYyJs7TpjpAfT4W13zmlx3G0C
7JhoAOPkAfchZQzi9pvDqei8ihBtu8iQCuGSC+LT04I8Rv3VHzxt+IkoOAzM
Nzl5yQrnSTJvAiiGYB6lmG+Dw0yvcUOA81EoffgYWogp5EibLNKDO+ekGZwF
1SYrPBG96bBm1yq/Gr7g3rYKdkBiUz5K7Jf5Ok7oPhIdHKPDBNG7dxOfWO7a
8XIbThx10wvuZbj2Yelcdj7gF6DVAidaJ7U1c6x6sffae7121FDorf9EWKHa
3B3vfH3ojhhIHpblXbq1TRJOsIgMTv62SZ6bHoItUV0rg6lvw1L8VPzMnliE
RIAQY1W2FBjEjaqv6+sMRJNTloPB/mLvPBN0/NXfTFkXS/Ga8VS9zGBwKJrj
tEwnmFflgIYTHGnSP2yNw990qnSJU39yM/uI1ESb+FF2VYFs60nTTZ+XaFhS
/aPZEuWOlP/sYq8PfW0fA6IiMhcN3SafXY6qAX3iI0q3b8zH2Y35ElUygUlw
YLe2CqRtFISu13JgUGXdB1m5GxioAdjOLVHZ4bIHScuRZ7bTA4X1H26q56EB
MmzqYEIm57EY3EynkbVMs9p2DICRnTOuOO3Eu0iD/vsH6ifKSHySQvFIRgtH
s3EbfkEhjTCXDq1dt5D4wbokBV/R37o2VhaIlg/eVM6zV9mrYU3Qf2uaw7iP
7j+oF9hKxHanCHtPac9JZy63Wq79UxJPP6t3g8s9qW4nCGcedkj65LWkRgjz
53gAP/ERy/LW/l1YffkzqYtPAIqimqHtGYos1vTtuZNHh/BXVEvbPGDj7jrM
aARIbp6xpzgff92DuWWpk0LmZe6sNOHJ85dc8WpxXsJPsuie9RbXnTd8lCdS
iQQZaO1USJH82DLClLlHkS4kJKuaDjC4aSrf3/VfTazXdgyeSFNuSahStPJL
VH2EZGIRFyGiihS30bo13aDbYOKDX+VDOQUxzYTgaMwrAcSAnOMTqGPRp5ON
CJlGoxl9m2X8uUfFCtCxSSg53K3S7RxhUPk0BKkjerbBSfBM+Ie4MpAG2uL5
rh4Ft1rXXHS5OJZ0k+TKLlFIJu4YqVUj+YKo3+lmhvVa/ZQO5l9UT1joRZqR
KcZe3dI7wvM+fQPPMUPd/kI02A2bYN3rz1LeD+q/Dk7N5gpnFUNuYCc3l/xr
qJKWdL712LAstR20xOrj/iLEAdJBcji6sheT8EU2uFy7jzPYZvVR40aMvP2S
CODgD9XODTkftk9ffOlnTXZok4jY/BDvnRgEWLu98tmtpNQRhWEd8AvaJp6W
AhYjTPXcrqDdX24/R2P7Mg4oPQHPKp8JnkrgBS6mNIT+2/7Vop6/2th2iVa6
KSDWsJEMgJtU/n/NVXX25scMEDjh9qTYEGF+Cg9G0BErhDCUsJ6Rf8PUkfSS
nOOQBD/tHimVIJ/FX9Zw06tivx1teOJfNaGg0PKGxbX4HFyM1mj4Ql8u/q+e
ugIXjdQzPH8wIK5eAZpAHl7qmt+R6Rr9GEI14/AEhigIhEL0ncegYJ/9YddR
k2HKltuL7sMgUuL93rPPtyd0tv3Ui9ep0APeAmn1UWSNm2FnWIWHhSlsv3rN
aBE7ZKdW/VmeiLi5fWsr9GW/RUqPKBSI8+IRdD6p78aBAvQJO3IsenURxlf6
L0MJNHTC7QHIkBArVTuMvua+2eULTxb7/8YibXeIp4cQPdDqEv0ZIt84BsBl
/UPPhimkb74GJPqfhKHSSTSTtVxKnGJzRY2o1EqOI+GhJuuES2+dS6FgfmYU
MGiyiWj9NjpSXIN6+Bmsutz4Fj4e2o3K9MThNtqy26WuNclSQj5hTokvDbP3
JZV38rCmHai731KTkbEuj4Ef9rAqTgKKosMT0/aZJmm9zLpNvBZhY5arJeGk
/Glq1KV83VjDTaaFevtnVdIp3Wl5PxRVEF5TqG8+YllQD8DFKxr9xlR7uG7J
X/yYNBewI1d8+JTzh4KLgYZisYol3OFWf6BJf/c+PjSJPL+SHYMHmHqFqnUW
HPUQ5wU0SAOV/jycgWFime6h5OWNGjtZ5I9t1W0ani2o9HjVwwBoIpZ2/wll
NcvIzALWrv+vIoIE4s1KDPL6oMvJnDaVUfahngEqTlwGZq+tQgxy0JmdmkPS
jprOF1TNYhuvcZPPQTmcye3f9IrKQP4dKO3QzGYpVm/ge2jmEO01GgPPFNGC
+fBPlRMzrbUMS4GmHYNM5SxorU9xuZcN2BW5dOJJGaX0Cl5SdZCl+Ls64uQi
L5XfR7+QdAJTUk95k1IvUN49zGgvJI5ar58Lyex8XU35aLfmojWzfPlnm8U0
XExs0csFOX3ViDol0PZAOu7SkYeGvC3l9oG6MJlWQDvqnOU81aB2/eiw5iNP
h1J7cyeNiSs/4PtgBHCehJTd58iunc6anQdqZjM28rhii1OczgKOF1AyKBeB
YKlUH8lZhiEXbaRZF7rHqZSpMq+iQa9DZvHW9aq2sH5v6SI9t6EunH3UKpWT
B9rB6QdMGBUprNghtmECmmIWpqpfIdguKXjloPMSpADdiZ6C7J16xqxb/b1f
pPIJ6Kfer0a/14eZ+3x40i0Vlqs/TsilltGe0Pzjaxz7BVaLg8STYPI43MvI
vboJJpSGr8GaZ9NtuI+7MDW2u0VW4Pt/lxLuaDbzAMwfVLrf3XbWGW9RlA3X
SIvkvxE2YHl37MNxHZOd+tTQV39PfS47j2bJhejirHW6Erj6i8sFnyOZ9I05
U85y74GDX7oz6sPJxszDnFSm7ygpZm4CIo5VAtc3PIDFMq0oVj/DCToMcuIC
YyZ+E2Iz0dH9FzPoH1q/2jFh/IdKgReR/gk4zhf0NzDbGhMuA7yaG0AHHPQQ
fowTBD4MCbpWoe9x3vcTnisRjSXDjWoFSQWONCGYZpmzibtju2Z5bd+g6Ics
1w1z9EooWdMy+3wL0aRJRcDEMciFIPcwQ+GWM560CkFP3B/910+RDGhdK9Xa
4z7s+tC1YjJFasQKZZwXRPVY1kOrXwpEdpJpswMJqVkUgakdnf6iSRlY6f24
0wcnrQhUAxlRTihLDsEb1ZXgza6XE9R6FBLxYdh+3ShPzjmI+nqQQYUwAnwv
/d7SaKvzrXcS2cGRydPHvtdSEEYv6bO1fPwi/zn0aWiewAHi0w0fcCzbExdy
B5dVoaPtB4nnZyU9amNEYjDMi8Om38pr9N+Wl/nvwTz1pqd7+h3R7oGJf0S6
rWFP2evHVnQZ9you++ItNamthOTausc+s9uW82RotTG8U1SeKCTLOtKN/xhZ
/gzkkOiGkJCUvoAz9ceWI1cHQsxh9KUhV8Zclzi66o2Ee58DCGEXJC5ZmrqV
L/nH4c6xiSdxCBsV5Tauv1iDWVqnRSr/VLi0/3jNsfvdYXEUUK6NN0hTyorg
kl4GKfjPBz90dKlK6WKxxHUxuScoad3qX8v0cLYNjsrj8ejRrerj0T5xAOTB
r4EQqX/E6YZmCPou8rgG1Q/EV9TftWGJ6hXcWMHeA5TMgGIP57VS2e8Jlz71
kcTv6aMn8ybC1EwEWAR1w9norLQCNtsT66dNfoPCoJsMt4n6ACVeyVqwmIGt
/9BsjicQmu4UoyrId8P1IJkH7LT09idMMxgJijNQIAJWhGGqD3wKyp0sFbDH
cGKggOgFc8o1CwMWSEloLk2op7J+gpDnVE/bMoaLSm1yohBeV64Q/hFr3q6j
mQ1FH/AEcQ8Ujst7zN+9dEMGvTynQTyC0qi9RWidcRqtpZ0djmIKKr7a+6ZB
kEsgJmbMPAa6JiyTQJHVzqbO5n4zTp7VbMBHUFyvoqV2PCYmQRAjviAlr3Hm
fcNtGfL1ylxG2PL/ptvWHA8nIMLYUUHU41HtdOfBiF1gkXPx1N5e1QUmJdiv
Ls9hcIzwg3TOw2Rr01nwPlKgGwSSnKKbu8hgGq/TNv6cPf+pEeUdIC2eynbZ
71OE3MNeM/4lhYhqdxMa+7oPPrCrHeLwy7eRScXYRAi/H7S2VpdUMZWojLvw
wer42QPPewYCTkPVSbuabWxzdEMPajm2Yu7CsAyNvXJvqyDpEcE4ud6BuCJ8
PGJeMv3kJu2Irbg3tEoU63LIXdl/Wg+WfelcT2z9BodHw9A6aMXGH4eMOEl2
l1xHX458PYiUjyZ4cAjtPonCuVs0W1RmSyvlz/1gH0DV+ThzJPeM1z7kfFVs
BZAcp4onBezG9TirZLBYjo3ixhfyAWHb8JKdMN7GQJPXrz1ek/3KhzhDfZ+S
7VHMaF8u2aWyJR9ZI9xmNcuHR4Fh+RdpBWYg+swSAMfpTRb/pKo5fjHsbS45
H61/6+lPsZqjFwSG6cDQB1h3aDkdcaQwuPsWu7TTz8jgdEU7PTkNZBmhZN02
Ov4Q/RpGx5udIOszdfhslWlsLR8R42KVh7ei/yWUZN76ewata2+Mh9cG/DDz
Z27QS7qmuYrl69yJl0LAGcMVhabnVfBKr4fUGkGpzRE7H9QtByFQcSD6rt7z
CmtMvwFOFo5FRs1kv9Gn2+8Yd9zs7bCjLY/3+E3La7fMgzpts7zqgzW7Zzn7
ymjdNpdVsrAOar8Gdo85vqPgwkj+2KxsguX32QTzd/fNv0LtSjFc3aDF8uQh
Gn3+zWKtJRV1kwWyYBU+Y49Jv86N/DCwK+oYTD/25dk1enanaOxt6cuVQ8og
PEMK0PqqWkZ7ryOZFiQcXjKH/L0FJo0UFcRi+ZwL0yRvTokXJOhkyoD45TvZ
UZIUmS2O2IvawNBD8IYPToGW2PrOH6moUJtb5jjvv+JUZFLu0r3RqntT4f1B
na7pewe8MfMaDHGjxf50Q0ARpC+s15Kh3kl6YhRVSC2JX4RW6wq3BvgxpLso
AYSOUMRQ3PcWuLCr1//75Ro0BkCXFZ6W7c6AXOzYiUjML5uPyuptoFvX2FZ8
X1sI3hU17Wtq3kMfWkfeQ63ETbilw16ZmFezlbtvLAW9GPaZBc3mfADl9DpY
TNjbUQLBHXPXGzGN3p68Rp9edPURoD4ReVMLcykhHu/60UR3lLNaNMgSdHqP
2utlQZH9Y1uol0UIcZjxExTerLhVicrP7ubIGlagzP5t+C+cLoho69+BB5n7
Qwgm5gFrFvtOAF1gC6v7/Pq5wfS1DkuRwejrQNbMyIcK7C0ntJ0swHlvww8T
uek/5aoER/S+Tr8P+o68/RVSpvk4JvvMiGuR6q9HccuaUSutJvIlEK0Txk5Y
jQBaKxxo03QVdturWLYAUzbdQYqEZwTFkm94AYp8BT6AOBDZrPqipbIu4tDG
PJltfiFF5ENz+96y12PqHNMRV1bN8s+YFD+lOnEtCT073xy/Tx+HOoG+ve+/
J1IGhi4UEKfW0kDP4ZjYuyiCC1Ta6MqXJ/75YSCODlZiDCC9mKH44gQC1Yh8
6NSBbNcXHmqV5vZEEWyKBL6WafeRLds3Qvjou/7XH1nuAzZWdHt/rt1xUp15
0CsrkCBBIlDZcRdkJuvn7vM2VWnJt5vJiMs3B29QDZ+ybZkOF1cJB7IAZieK
6B2XsnUsFquZ0f7xinUmDLWn7rfqWPRuuFYZpypzQnmHP23GfWP29bpjOkar
kLrr6iUTc4Xcw8jH9DMrfEQZ/4Jjzhg8tAcFR9PCVFTXWdvPbM8o5hWZ88mn
KsToZX/zXwgKSeUlzEdtMhjzx+7hko1jOPvmhF42LoXYe6feEu9JgZddAtjB
ngiI4BcxyJyPv4DrC/sm0HfxHi5mbpfrHnN06WMHScncesTwXirZt2Ml7zv/
cuuaqZrEjSPxj+vgdptTd6rL9KqJ5OdgK5mX4jAXt7oAt0QM4+8zkt9qxswY
QWW3QvGl0YPiPHvAtUjvOvojMezxRyS8dUmEsMtHMh28OEvZ0x9KZJ5xgBde
nPD4EESjquyJCDcGZsS6rn2XZMadg1IBGhH092JG7P3x3BIcMeDpvR2pIi3k
i+sBsVueQisAfxAOtjw75DpcVgjfROWrx1em1p8JWiOeMxFlRswWM9Es7h4T
ujV1g3BtqbTzrWFM1xydRuCH7f4cdQdiyJOiVTEoUiaDs0aQkqzC9a1ZCLlj
EDC9/UHcwjAQTehrZmTnH0UJeizYBUV8X7Xadz63umMzb0cWg1t2g0IZd3L7
mRXQKdhM4mKD1oYH8I+4uMYGZ4veROxLIpoCV6JZgd6fuNoJ4smiGT/piZwH
KhWx7OkHZafpmi4HSQmelzTSI+Z/pR0bxEflMdYQKEIrxP1R+0vWNBKxpU5Z
KG7YgiUj84fnTuookvWdr0ePmIzDjHMDmvCSj/GS42/ShH932fsys2BePScI
0d8b/6DJuEeAKviLSPovKW4pzkP64MCVoU0K/Nn4NG8x+ZqPWmbMAUcHch/5
O9AFJ7w8ph04ibnLcpEpogKPfcyocMGhStU9RaB9S2cKkYtNl7/NWJc005ay
QdCaZgokuPrYhyoFlOw4Bj1WufBmfOPkXaiH+9giIp74cSjM9yBkWFsJyHsr
gxkjO+RRosia1KhzMyFpomF5Bcl3kxvGiA2k2Jp2Xj2p7gLa787w3PGzaOgV
ySfaNbpK71FSJcksIaks9Tn9M93bcshDrAb3hmAnqG9ivc5ntaZfdvQ/sicC
nXU53NrqKleismz4y3QR4JT6O+06MCXgp7vsQg70Y5yZ5KVwPTivwEmfaETa
YK/alW9D+VjVMz22vEc9RQISnpdMsLkGFfweoV/JaJIzdvoBPkQfrGfDv1O/
Mu2yoSZdN1FGuxGiwmUsyfBGX50QbZrSjtShZ1th1cIjHqDUhrF5gqDlvgJZ
nOLApX2rpUgi7jhnWnnTaXvjmUS0MnLqVA+cdU0L67ambRQhMwtpdJU22Ze8
/jTniFdvYBHoASMR9ZXeIoCTOJOtnUk4KecHHBq2RvHZtEAWR1sjaoNFbvdQ
RbeRmFRxjA3xECLJeh58bpjTthnTzWn9UjQtu4KpVi9zdVWul63AKNwHbhrj
aTGDiqoyxU3ktu7weezv6ngX3C6tR5Gtg9b5OcvWQWudpDtzIcqtdE2uNz97
1pKcoUfwfp3LjXR5B+mWhV1YPGTUrav9DU/Z6ylx8/GL6weOrlMQQL3OJsrf
3LeG6oiclhpqK06954wutEf1Myv6lqsO9a5+TVxfyEdIzbzynsFH/0K1okG4
uO7yX29lO0HL4LQ9sc5MRQmbLaJk25qrwRpFQMD/d0BJx2UwHOAsAyTjq56f
sV/XDsuPq7CqAH8Tq1SHVsibkztA/DOriq74/4K4xNBpBwyx/EuHqZZHAdiQ
YyFvO0LAO6CpyxH0GYVCie8AiOq7suFkaL4EkxCkivC9AJ/2U37ZTioZxhCJ
/WQyQIji0MQFjvXBFZhgbuT3Pf6wk/TFiqxjtPlwi6VodHczNexq8JYgxIu7
U0tZD4K7BAeJ+OKzKdtUyXxxi5RBgrzF6hM+WavdcQFn7BLfdXJ2Am5KIm5W
Ix45Lk/eKSfcjskYHfIZvU+wwhGONwaBg6kCwzpAb07dq7z4RafJFom1jSvg
aTLBilmEKR5nQWv0RAgBlyZ1z0YQjL9D2oUViAi6Lrx/1BqpL8sAZnBnJ6Ir
JHo9i5rdsC4PzOMR8W2K48ghTClniWI3rzjIPb53RPsNdEseNXCcb+bfDmUF
ntDyK2MKn0nAM/lyok7cUnZI8TgnRYrU8pYlFHcA1OaNNRriyERu6mVvZz+K
ePr4k9BsH1QHFo4xrz6cddIGsGnftFyB44ASK++Xx5OkZUu+G/iFecolBvbH
uNUAM9GUiteYcDhFaBAGCw21EX7YqZWng9XAWx0KwIlzc5NKzcFSbaRISa7k
O1tjzubvyMcIWiQcD8xnVtQPhZaIh8GsQu8izm3Q3v1wVjktz0neVFLtTh7S
Y4wXfTQj3jiW+3razDFhTpjGiK38vJ3PLpYCkFdAJ37as3CkpbFBiyt2KS5L
7jYMYN72nOBqZTgJpCGvnNonyyRbkbfuvSRc7zxZJdSb0huMTO7ZePOXCgYl
6p/z2COiwm7Io0J9xkppVLF2gRMkjX77g2IXHfLX4psjocYS67xAXPc2NLrj
W5gmtkMwJinwJ0/wQklkf1PrwebRw17hSW3ZnKfHZdFvwT0GhVlPZliXSyZ3
yVuX/lkwM4xLdkcsdUi7AteAF7tFkmthB+WEn7BdYE+Gvmt7oKC0pKbIKGvW
5raUGICMsJ3fO+i/J45le6wiyKgZk045f3kD6Y1W6z9JSVDng+BDlR1Y9ffb
nnvvS5/gS4K+tlUHikBTdfQz9OKQMZSqGC2MC1FkymXjKH7v4R5L6X9tSdsu
iQ89an/QicAXJanrsko0MN7uXNuUwTfpY99ODTmWeJ2xcNUHIpJRHQVlykV2
CmrC3lGnsZDCxn0xfo7TIFsRbGHW3UCE1+xj1LLSiSrCXuihFCE7n/CYYowE
wNkWPzk8x5fh3LNYozaYcywH6jJyHfILa5A4kYQoUBiugB2I3AwljOxGeiMN
YJU+v+POhF7Qlwf+HZklO/gaqmWbocglbIJuHobKdcVaGAcdLjmN8nXybrey
nS1v3zM5/KyMiaRXNxsh1xU/KBc8fuUCd4FRyZLRbFLHS79L5ZcZsucK+Qa/
uiVRJMsXpXkgXfRAf+lykh8keLlG5fIbtAj/1UVIlRvzGC8I5KHFwX1bB3w1
L2eEmhv9w/e7ZxtoXLVsB4xNsHcbQxPGp9dlEVC1a63SBaIQqmXfmnZ6m9pz
hyNfhh8wNFwx1dEdlpKT9x/X+GLmWcDvlo2ql+1ULQ9sbgMwMniDNzA/2XZ0
7pGkvS0/RiDQe5bv+LFk7lfj8MYoN85z3p5vmSRwyzO6usOPWu10oRcvYOAk
L/ar1YhLroUpZHR1A3Z9lZicfQ0+16QU4Ggbc2ERZx2qttYA48/QSlmgbHEF
Hmk88bQmpDtBreQSQ2nvlnlkfXnt3qi0H39MfJKINWfE7s0nnBl3P8QOK4at
EBybBX7SXCZRytE1XPMRd/BCy4SmM5eape7TsnI8yPu8JsqNmAaYbve+MVp8
L2KMRtpSKkyuDJ91xdnrrh+15+PDoxmlBDJRvfUE8pi1/vH3pEpQx+tS40d5
LjPPHmeM+68xsYiyKraAo7eK+spGzkvdo8s8rGMdT4JWdPWaRHD3zjgimC8D
RJUBM7GhjViN84PqU97P9VAXJbail0pCBuJBZbE6z2J2nEpBHDuotL2soM+1
rBIuk4yABCI0iPmTS3GPn5Eb3osxQTdTtaVkmGYN9PHz+JLSvdWNms53tO6s
B76n7zqCpp0WoiFSefF4H3reIB+OuHIjABpvUjUNiYGbsJswHmExTPr5PGMM
cSL4BOcMC4kaxnnLyUtzwJZxlG0RtBPPCuH6e20Ef3Fv2CdOgEjXp27BJAb3
eZoyIfH8COOwzFcTypcb6lknXU26RWZZ/jKrrsCdIqw4RqZpi5csSf8N6bIO
gO0FX09J5FS34pJji4i2EpPfEN76vsvLnWDAjX/pMKCSUfQAzDUMcZk8l+9G
Ylx+tfleAeOQ9NnXoJsBPfJY4493DAEtVNj2jDQ0uHd/tLePKpqV9c3HsOnp
IyB2m1LJDnzs7SlmKv7jtBDfUeAo/zfNZSDZuoWwMCvoS1bI/z+5YI9WYHn+
jzLaKBmWcuQHtlF8neRGR9nGiZfAXtRXLIPm0V6zC6mi8+HVdDouk48V/mkS
eV2eZaBKiT7c/aHujsIPxk1UAYhu8mMjwTQJRsnFHTO+7evLAQ7TqKgU2p/G
rpkBB8Z1inT77y6HGX2iOYRSgc8PLeLculsvTHu2Y6TVha3pPteEnZcHIjs5
N41zABUuv9ccVTZIdTOLsvhLEvCJiIdWs5jU8/CbAE9UFwFGrjkLMhDhdm0L
yaNGdzbX5TQX20QO6uvKop9eCnIdKg87aVJ2/eXMh8JSng6jBesDr9xvLQFN
HZfsNvRz6aSrqD780TJpVe3jXMWwbstEQbGgFztoyKWEedKWvJCa8wYSpjNQ
l3g4ahQ4wWpSL33mqKDOCb1RXppdrVyk85UPH1x7g+YlSzTiw5MqAZliuVTW
FhHC3W9IPwyqxPVvCY+HbyIE8mYw+A9aEOWerF6PF7cN4Nhy7YlhJ2Q3lQOe
VIyTr/r5QI4ELzicXYaugsnj4YBb7dKkilHiM8Uy77FRNDRxnhJKYXzp+DGT
2n3f1pywQcMU32GYVyF8oahhK+z+TGNUnuUNS87jML8AneVyF1uvnt9HYdQx
sORKFcsi3hTkRPovcJDKzGE+SlQ9elqGLNBXctnX+MpLiOHud2FbW3JiSYQ9
/T2JOWHZtn9JSbn22gefSXqrUk7mKRaeqTjgCoZMZ9hkf8j/tWthgozKUyf9
omkFUrCeqK6nnOOi+lj9vNpZ642UG2jH5OncorpCUaudnjqygz7HDUE14YkF
EBj38+sJCOkyxH5t1HqBP4VTPG4BjDcVC+3D6gBOzxWjZcX5k9sQOJ13z1oj
djbxe0flwoKDl6PY8i19r1fEYc2w4qZPbhn69Aq+PFoHtNJFgeL/dXyxVO+h
nyhJlcHCUKuzd7zrp/BUz5AqlRsjpaMK2RtYio83gXlbZYXHSRbgoB7+WIQ4
FORaDhpoYHMsEqKgWO3BP/dVxt24GDJ5Wz02+f+HwTwMd81El1GaNL8Fkyjd
51pP3PwkbUaHSAZvAQvxeyaDNSaWaC1llIO2VF9kSv4MyoxSzPZ5qp5bljSE
1FyG5KwFb7KbMHcUWvfAsw/ZP7n5m0DoN6Vrao1N0nA9f8htKxhxxSr6x/+k
gqBXnXKkS+oi9tlMrpJn69hqe29rsu1JlthnFXRQkkgyUvHzMauq17NA5Rt4
DZVCSsm+KxcqYBEVHGL4My+UWzettQBf37Qe3l3R97sukYmT1Jy2qqnMz0yM
OjTwZyDK0Sbvxf449MZk22pSYMvJ18CoBMUNyV0beeVe1W0OsvXglg39G/GJ
CK64MjRQN3V04BDrLrETLrRZ47TUJ40DVbpIuD0WiB5jWsDFpW4j9RNCc/4V
+vauW8wzmGZF2J7yReBt2pttLBbva6QRpDQsiV6cQ1jvaUNUXCwvo9pfMNCF
/cUIXAlpZQA9bvZz9RuBe2DeJOUSJVf6846tcpvVc8Ee+5YX5tbnkJsa7Prr
hbIQlSms4GPKQWS3CCvoJ4TQZjqFRxY/u/mj1bDMyqi4k1HdJR/EWBv6tBeQ
pfBleZZEfSo1GeXH/k6RtlAxkKsOlQbSejvG+FbuwZ2lxH5NxM1l7zuPRj5A
GLMr/zeS8LWGbem7L7Dnqhhm9XK8Yn0sgj4vUj+k+TqT5hoRpfpOjM+S+Ssm
R1bQ1Nu/YWIGFo4MrryzxditFnIxIjBp9q241dW10anj7sPDq7nOt3L8rWGJ
o2mMSdQl7jgyGqGheAwRX+kvlg3j+2VGRlm3xmAr3ida/jErnjj2faTXGuC6
E9ylPAnBhzT7ZuZ8EQ7O4KxKM87N9VpbuizTyykb910NcS4XfSjYY+hBXSxi
bq9FsQMhB0uZmPeXAghEE7ya03Qh207dOANuLvkLKFKxRW5S/v6dXrzXuhHt
nAPaYSC4suk2TBrVickzKLjQI5U1u+xmOFBE9rAbaAQbvBM+jOPS5iiDEu6r
mtTpNDUsE2T/rkIi41PzWu9iEz6CuH2bB7RU6Og8CSxgxStVSfnUEGORZkNn
Q/1e61AMu8nS6QJl3Jb3DtyhKkp48KeLYgUbhLv/yKGgDdqK1MT2Fp9CoZEa
A8mSGe/whF/ajwMbEcLeHJQrO08tQZsOER6cZjPyqMKHkrnTAkOwsLS58MQT
52226Mchete6kWaKau4WRyTR6LYWDGI5Zdcz6alf/WNFoPIb7N/AfObfYTNH
HXeeIWZ1W7sMf71Zd/3oCSfd9cN545v5qXOFmfUImuTqYurRmTjsMyyCFrC8
GWLQ5pGToR9ldHMMcNam3sdbfMXOMcXmExu4gC2onZpsycPmvjaRGjJYqA5L
f3yKLQ2bLRzZUeONwBkZA6SYKvcJgdNXSV3q4rTYGL6VCqEKrM5vVj7F8For
cWwa3yo9kTC/570QlB/Ri0Y2v+h/0CUC5OyKHknvZezRw/nvgCeXAtulwrEZ
ttYXEMa0BszYrg8weSv1bmA8PiUM3x6GG19Zw/s4+V9vAgYGEPekrNtmwvi/
ivBCeG4tT50JzVNYYZCBAn217f8HawMGU9F0JAqq08JM73PbIt7PSaQFIKJ2
s8/y/88SGubGA1LHjucyD/VJzC6LnmeDSZ6vgjbTGl1PF8kii+zmN1PT5EJ3
lk5L/AkJxKwWzxpD2XuJH3lGv4W31v93m82CxUUwIJMmaMCpilHifs+b/ryd
UMW0wRqHzht7xD8qHYh9x9w/T5TxSQrsoP/kper+Ls5XzsmzFtBu4J+jHdR1
4lB4R96FJwFJycT3OQ54gBMlOtHMU7seq3KeoOnl2cLyu7C5vEX3u9IPOZqZ
YDcj4CG1nz40oEeXSMGtu4937Z7g3UsLBNw7VZjZ2ur/Z20O1mV486rykj2b
Yp8Eyjg/NZ5uVifCG4hMaRwv95nwvcVXFj64OXnj4X7CHG1q2TRmSoLDvc0Z
xs4tzawTD+jAjrW/M50BMbxjGliGiKi/9dIy8/cE8nqrvEH4537nkuEv0K2S
IR4QKPrCWuOo/hfzebs1kOQ+JxLB1cdnl6gPvw7NoejM0+rzRuzaoLlQqQED
FzTBFc/BlrywL/WRq+6HwjTIWUMm0UEySiCGFpF1gVbW+ftvkG0YjtEIVXXn
OJQf188wFOj9MqEUpYhMCAM3/uUT9ZYij/f2G3lvB72NXUFV6YfCYgJ4kMxd
Zt+S8rfu55ZvrMF1PqQ4+vy3k2dZAlbBlOlyTrEFzy5B5+vbyo/q261kczMM
7CpghC0bPNYhhwOq84WoFYETIkPydHe2QBxFeyftClqda/sGGxzSS4/baPIu
XLE+qXHg0NoC7R6fI8nX29/Sbit0EYUKXv30CWmXuCXWmfC1zB8kdFDm5p/E
F8zCX2IHrzjcK7W1qbgHd8rUzd48rN1xjdxA/taiO4jNKbjd0wtH1cwtA6st
3eKwvx1R5roKfx33fs5V0duuK3fbsddTTSCch1WvQlUgN57faHR11EpKFYUa
RTcwmsW9kKyAFTR25a4jDxQIP9V3eFl1yEg2vsqyDC41GATBuG9WbWfY8auf
exdxRf0uKEWx6j7hHQP/R1kz+bHtrkotnZ238a7V2/Z+KcSetCxV70YdIdl6
9JR4YbBFcSKuniJcM8LnyEd4lb6TwWHhg3KW7zg3YGpyjTAUFWHA2EJf5geP
kukw5OZvZ2gJo1Z+B7FaYeVlHAa7+tqgzs3H6oJJi2rzDp9Th537XU/WbxA6
qLJFNL2K0BU9TTjDOQOx2UFX/Ob3elsOXKH0qAR4YXoLmDMEV9UBNQ9B0yvN
EVWbXQ3ZQ+ljwgxULhORcxWYJhNfkTbXYd5x+hA8nFDG4wIFie5Hfy/75xvz
jKIhQgQDSTgW4Rfva4Xq61U8tLg7Uqk57fjQxXhdRI5MBJUp1dauPlk8fPLl
pgsoFPYjNr6q8T6pCdhMHaWxrQiEvYX7C0MJ89NlMfqC7FBxV4CAMq9CnGzC
k39FSfErdOuhbl8PJdobvI/P49EX3LL9x/kp+Bo0B5TrWN/QyuEsoWeSZjuE
835dxLDJstM2W35fhkEijanOCcJDgKkUKxkIuT/CV/VXehwwj9WHcwl68z+7
h12nQ+Ce9kqArIxxu05GHW5KMJjaIN1h+gY88xX9mpyUv1lwaaXYFEGENiwK
lW2VZKh+Q7b6kQSQkHLrCr9aBJa7ZUtp4jlrtT+d/N8sDSfkZDIZ41W0nG6H
aKGn7G2n4NAR6A56HygAuswbZmhB0IpMxUms+O/p3FYXr+GyFWPSdNo7YBKG
tvuJqsuSHMjaEGQ91tpVaPE3bLSJLw1TXvCEHUTT9dsQgjHqJ5zOuxcfbVwf
eEjpw5Eq6eybCAeP10g6zm9eh0amyvwjxKrT+OB+2vCyQFp/6YJtmdsVPe0u
+aZvSUsw0PFzMzOiEQw4Zt/vhUc1qIL+20pqju6Utc739rhvmQedE+59zP/7
fTfg30sWrQjf5c1IwQCwX/1xBmnFKjt4go56Ulsv1tpspR3ZZtDTd1abS8QH
ByzLfGmB9bNFVeQEDlwYFzgEqhbGFIbkrdhZNActbc6lgof5xHe8aHZoHwNM
9HVOuheZOMWVOLpWWiSvMKMpgEl1upTB4lCaJj6GsQFaRDPp5caB6kP3C2W8
ng13kqhplt0g8v2RH/Ax4/rht6gek/S9Fv6W1l/fi296iEZBNCUidBOglXnl
4ICW8FFhHXHyJ4vjfrqlxsB531mOatn/HPuX2keButvBITaKH0NJoYLEO4jw
D+JfUZKydrDkFoPcxt3YX9hJbk6ZB3kOIQksOvvZRwVh1WTzm2eG9rpmVEFS
eSc9QuVNla3ETuQSxH4eb/cggJExtawUC1xNLyC7Ot2ZZUCq9eXUEmBhorYl
JqUkD6I3+KAlIqTfN2uBfHTumLvYcADz16ryucsWAZvm6X3Cp3KHh/Nrvnqj
LKugOf0D3A8gev8h/e+vfvuEVwSxzaqTh96BQPE79zOzad5utEnEgi72AqSa
TeKAKwDATkHo17ki9edP+RbD0Fm6SIh1/VFwbRQzoIdyyqlxGaX7CitwKSH8
DkofZKtkZT7F8OpUMn2sqIb/OADcXMpAUfdLwghbDyT5zb4AG6R60YLU09q7
p485nfjdd9H3V+Rsl+FVzvroYxlKz9sdKZ2UkRpoExfsjlegrNUfktTQFfRv
4BS2nkymNvDmuPWaS8wotjr28p2vhafFdUGHcfYqhwcylsDDnik97P1j8qht
4pbCFHmNeWrZilIpWYEuwyxBjw8VAZD2kP0vjf8pvCqG5vfa0bXUz2K9MI2w
slY7ZxTpUfGBB8bBuTWWe1KGIIRdfWXiLV6trW6tdf3ISgv1Xpixq96N5zEx
EEU7pA10JBxuC6an4eQXpJM8ZYFk09zRnOudhRrJ96dYxzxtL5ASg2Nywr8D
kfw3mq6LQeFDYSAgfhBTXCplGUDtKUHtormK+FyD26clq/7Ijvi/bZKSDjN+
wmstkYSyXGqgTBC+iE1zJhvhBbjiKKhzPudxmjaEazitRDS//MXoXM+Q1ESi
4HOK8YmoUYXkhFUegy54EUYWHCjas43dBj5D+OcrrGqvkSe+7bHcq1Q9AkOP
MW+NAwV+9c95pvZHW40MHiYMmwmZQ8Rpodj8BUsuFbs2FcJRqZSa+dnHIKkf
KZ9Xq2WHCLxzcvKffSR9BxJhXEbFcKGuhnY0oJ14+kBJzsxpxPTMoacDSQNP
epWAN3pv0qkAPTJumotvCbSA7jcXoGpB4v285KJs4qcSGphUZn/aNtQElwat
tez15jTZ8c3V8jiyoJQl+EgYZ/RUQDJEZj9OnMz2fnrMnzaV5T91Pi2znJnM
oLtG1ezII9GGTZKpdrkXyO0IWJv9FHWgWiGmRsgEjcNcgFzChB8bzQVZi7Y8
H0kiuaHPvSpxVtoeckz0WGjd04+449URgwmBbqmDGCH24oNV3KEkIHdRp7Cf
nacHrl05gFgjA+vGZNrHHv8OJe3Q6AAU/w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI2IIjuhOXPPS6sXAXId2O9yrfexNLTLimnouAL4btoKfwOQ8Ctc+ka0efpbbZslmc/3NDQIl4f+jlgmQVDCkHFt/XGmUcYK97B+xUjUgd8CliIVI2aVs7mlSLK2kB2TKD0Q2q5UIioI2dimS6eQTdZh5IQLeiavyUCgRFxajg5WFlSQXqaHAYDV+//yHFWlVjipTiuPh2BA24DIUa889oswYsPiTbC9tm24d0mZ0dYr77EPjNydh39qLfrVgSKdZz0NJPgDEEpbjBzzekQ/V3h9xworQG36xXK/ySl3Qsy/zOZ9Aq9HUNUfIMonLIcE13Mm86DkDiQmFB+DRT1DsL/Jqbwg3q8U/IpYzEe2Tghke7lL/nextF4NZxpb0yyP57mZCKskOdn+wa/GNrUWvRojOvPmoFNuX1X43tDJP8UhCOCIeJpf8RRyG3ceEOBaVyjhgvPkuaul8itCGKRu4q1cASt/r5LNFk9b5bsn/aIMnoDGyeGFfqoJ2iMHRUB6IGeDVRiGwOj3dOrI80R6foUGBuHSusT60RsoUuCfXK+71YFJ67C2MK1260hs2eKFt/xjsXrZcyx5L+XI2jiy22WraKIm0Tf9e0+Kv9OUEEbOxNbblDUww3bpY5VEJWVfqucNZjGAZMYmpyzqOSm/XnVyEHLu+b7V+Ipwz92p9xrGkaYA3vefG3Iz8qHnClUUjvv0CwHGM7rcN83tQj3B8RPjQDm7KrSwUmImGmBwbP02hYgru99bXYLjbNGF4c4IcH//VwmPk+UILcuDmehgBQps"
`endif
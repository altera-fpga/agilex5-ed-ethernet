//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MICP8fpAgbLyOxZJvmKK8lrcBuHAHDxSIf0RBmJxLdTaDHyooggs1a/zTiup
pBv4y8zlVe7fkz/p3M26IsRPJWtuHHJ6CkLdkNFpcSP5PMXC9flpp+76a+3o
0xHvPWb2WhL+GfY7r6N9Y/wsdkC34CQImMNV3eOvaeom03eX9k6uWgpqSJ3s
eVA4Ob/HJhPJTbvqD9P3ol/Y+XutxXLFYu5zJjcKWVMpIR61dpQk6AmgBQge
1FFRcQOffgrQEw6ZExWKXh1fRFtejNLuVW722zcOIIdgScLWrgsTrWiXuypf
EyxyruXH98vVhpr57sl+NNMG6+c1Mal9D/YCC7CnPA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IabvWGMNW95XMpWFXhLzlnOShawSyxrgprch2G3QD794+VG+NZEUUDYrdeKH
CpFaVBZtg7IKyg7h0XR/+DKHLOoiwLJpM2E0yEyROqCz1tqI4D7PU9amUX5v
zttQX3p3R1Ej/edAzqDe/qazbnH3Rnw4oyOYgvPYk5rRUhEIh2KR8NG8Neo1
6PmvQUM/Z31qC0G6X7LluSvOqfgEkzSLze3YEuyRMuPEfpFlXwwNGYwsP0aT
unJoseyO11AjHgZkYzcCtr3VbjocDYT+vZmE+ngY+R07xHdpr3jHCPhSZumt
D69zTwQWvBJjCX7g0H3qbRhksq9XU7Ho6m+iVlHrUQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JDc2YecAtGBxQLjySDzA5KGqhjFKr0aN1TmuuOBbsMNmtrlqcUbxU2TVX56c
GjPVvcBBCLj55RyKvQvjV7+7PZaxmOrA8FtTbB66xCv/7lRuhts/MjutmgUA
0XlVOKvpnnW0q9i7oRY/6/WRQe2HrztPoXVTBuLcz3BCf7lAWnb+dni+cCea
wtQ3QprUtATpckR+5LrHSsgbfkiV+qkhzsbBlcbPSd6y7dygUP1qc3dmDdKd
+hW6bEEbi/Z4E833IJqisP78HHQvwBvMgeFZcRn5uSEmIKFij3ynwUJNdQ7I
ljXYxgakZkUsjNvBzd0Gn4YkW5fPk/PV8YKabMae8A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OfV4jUAAIosJHDmtF9qSq208LIZUbmvkBHjeiOwmVDyWah17uTGgpmNmocht
OithjMedSUV0Di7IGxvj9qrtdqkUdZsWiHbJuiIxVlw8a3YEWLe/gc+Jg2jZ
Axvoy3B+5zrHmow1qipDzgfOye0xHxg/KnmXt+ObOwm9SiM6hDOmD8Ba0S5y
TZnmihD8csMJyAyfKO1rAhdj7yI4ISPP7VKlUpBZdxVMpN5TGLMlboW5Gvcx
EvkzL9L//A3ToMoZPVIYGh7ZEBBFrgNS3mRl3OZc1aOeU1KUDngARBrC8v5x
1/0UiRVBnuP9t5schpYy8NoAA5aIeOLvizqRah+tGw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qd8lkMN2jM9iM400Goax7EqwC0q4U8CqITHltAbr/9AxZ5+rSPmDaFw4qSAJ
BZ2Iiqw6bF7sFpsQnJrOXxXi574icfUxPRMFHJGc9lF/YHcGAQ1KVakR+fQI
D7FrXL7Edk3LLFc5aQC7d7VxpF2QeofrnQJVlj4BO3PNMMQhq9c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aOP/z3Xyq06TKg4nLLeOJY5gHfgCVqL2RBVum6u4epQwWmzKQTtE7z8uOkoe
Iwt52EtdsNFpIrGPmBIg40XYepclsSNPoxGQP/kob+mLFr31KfKl0pX5T47z
kBgZrARZ6u636UEFa3eKYrWC+VjJLyfGgSyYpR//RN5YdVM0HJLIDdEj8Kjm
aYtdpfYJHoiD5OClUW3Zeec8FScV5hJMi2oE4YTw79We6FknJOUjcSpQI5yr
1e+Kn+IuGJmZji63/3VhuY3RYiy8TWFnlrrv4rAChh0p9DznJf1nTpwc15Ox
XOAAUZSoWSUSPMRCv2M2iyLJfbctH9JN5P/AuagXeWFCdbfE0H9nPZ7vMDNg
gPvbzQl4LC0663p1GQYPmJ6r9pVbR5RTcvS6yg017N1SgJRTwqsErGf+elVe
uOGKYOg78MUhdxwZVZ1FfCYx8Pk6a8EtEiybVg8i4y6uMK9TQwUxGoY+uYAd
fM5AQXahhxipHHoM4JFtQpsz7n/vp/GQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
X12U4jGwvdYLBvhVu1XbOvgYUFlT/t/XdnjCA8TvMtfHMSO7ppbGPDAXP/Qk
oGMQBouWAdzlsHwlNtV4ABvfJd3NK1zqqitxtqNQ+IgPOrSIyO/sDQtR66SE
GnJQvDDJIhFewHr2LAY1I05Dm4vdL/LGEVGmvYlrjtTs9BuFGfM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NIPpg8xz14rdN+uKS3L8E41t8Fo8LHKex++nzjExcCLQKfrNwLoQgh+kqc0V
My0SsgbkMARaEqksYNk6qcJdei0rgTSgXLGeZlwZDZbx1AwYoaFIGOMgTY90
6M9IEEkcu6gIRKMh/nkl6O5NXDTuUB2jwhAGUBe4p+8cnKXjC7c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 64464)
`pragma protect data_block
+iCnq+EMn+34LdRShaJ6ABZBcbIBdiSI/Al478IxDFHtTdRkdTcAlotAReqT
+nlWC+Tkqd9SrLP8a9g+zw1ZWgqx3AXPl3+BuhjTkXOFMMBVXigeVpFQYEoD
ejf0nYsMGjRa80M3M+f4O0jIiT4roJ1Dl5QBgO/6wUCBjpwSVLGZc8zfmhWK
nBpFPOz7ex5MStuJyHope0Jyx31Tc/xqWCYXoSHHnjjaTXODaojgnPwfZYxy
Gjdt9/NOZoeSJjMFL3U93Hw7OLzULVkIFDHNbWqeKmVv0lyghNFz8+yA2dcG
C51FplQBheV5x9ykQCR4qiiVvyOQR3/vPw+HCO3t2qjWwmDhxXI2LjdJPG+E
jbgcHvchKi8PQIzjX2lRzsva1vO1BkZIhR8aqvfzzxcrYTSyfrs/2gLMSyyS
gfsrne3PoWrwXPuU38ZCMsJqLd1U/abj51etolA2yUizieuv0jsq/uq/0OjY
tvZZ4vaDCT2/sOTCvIv0wxyqMNtA03XLb3IjnAeHkPKPbuLQnIg66CF0tPHx
UZvFbZOOB9HFcx8eP6rtke5xkVyfVHtaOIm7vb1LbceWKTxNuwOiaYCgMIqE
/pwccU07LHUASCioupR6Rp6QD+ZnV0YgQk2SBlMS1J7niktZCoxI2XEbibxO
maJvs7bA+m93OaEUi169miBzWhIDRRiLIiTDR6RbTCx3thiI6HnI4luinwtS
No+EFAzpieGjYFwxmMVBCayhFa64q4AEL7eA/zvJ4a92HikAlYkPcI9W1QYF
YsXrzPmo5ZSd+Un1YOta8YXF6IvKEUf5GcpigpwFmblPdFz/gMcp1b67J0fG
VRUmvvDZrrrZHzsRJslXnhyKmG/37u7NGpvkuNaMxVvOfFiL5WkFwPf+eZzy
fh8VGQsMUFoR4N1vYgGt6nenueoXUTptGbLmpi26oc5qs8aIqYEtgoYxmF2E
k1AYaGOYnrxANsMFewKfPKGJLenLm3YCAQlKJwRJvcYNnrKkdsKaM4syOCof
3+itiKIUdlg+gYMl5Ene5KROzHfnUpZjOqmFQVo3NCMWJP6V2vAso7pSd6fc
DJ52HGtpT9dmKEo6FPK6rbW6zyZMLfrsYZPYudEF8JByLe1JyH9KbN/6O1Zd
nVgJ+tkmSh3XnX0I6blU1yRBizwtIW5wewcuI877K9l2l5+iRctaDAYoROMa
Vf9c80mIb1WlEG2Jj0lCOgzgA+JeyAIoZM6ql4aJC+H1U1/8baXZpRjcgSzr
Wcby2TgOdJsny7YYyg5iCSOcxlC6ikPlaqq60Ba3vcx4cEmuJuSR1FBaSIsH
WwSQbvlCMwftb7D5isONPA/GGhHR1iTTKr+vKRiCSashULS+Tj50J3mhikrW
hxgiRvQQQBzt6wFOZVlZxCzFbnYVALME4pazYwQ5sZTWdLSVvOLUsA2hW36X
TMz2qsU0EZbxb+TeXnMJMiKj6l/I0cIrCmtOJcqotsaUeAPMD5f/gGeCU3fb
pzQZbzJSFQVODbLcux838UySg2kriT+5wtLrTEucR0AsQeTKTj6CCtwbROmC
6uYuYE7sOrUNTam48sZYcy+fRWCPm07ngsN2U5134OqhyYSyX8IZOoTj7zPX
Nnk7pkbyCwhJ31swn4WDjk+KAyWSnNvSG3LkCm5aO4LKyj30Noyfsq5MJc9F
UUHUiM/u2ZoWNm2Ia6R3Mu5PPasKjcmkrh9zJ+WJPfpJWUjsqXGnUZcDsdpg
NWaZiVqAhQemEHLLe8a5z4008GDZIePKa+qg4gijT5V/U873CNd9/Chl/beB
Huf+gRXxmW6f56bejL3Ez1DJgwx93VbIQbCkpaJMVteqD868UE4141TXDRvs
Kw2ErhMt7sVBhRopOHMEwDV8FyHfT0xzFWBEiY6ewIv1b+0ScyjFEdJrXp7W
YqPJ/9QIdlTKS/wfjJuMRmLg+2j1FWKK001Jm/jfxak5p7F84t8P0VyI8CRR
8yagZFVzoLyjrWVLqyTsk6+DFAeQkfEAM/xPEEyjU9JmsoLvR8o5YW72fcaS
YSRrAj7QKAuCdMXrwjsbuOHrxfaWgTNKaYHeyvqRXwYg6NjyTPAcooB2zkw1
oZqGPfPStgbdSeBOGJ4VmcGpMe8DHr/7Doc1lkLfMUpbp616Y7xuUm3y9EP7
8Kr2kshMqnH5F1K7o0dk/J1H3X9N3AnvuQOmlypXmi/dabaSbHPZz7XyzUZb
hCimhjUMURKiCs/SuDo0VDS3ErFzShq5gh8DvWyGUHkBrPSfquq1kQhBy09b
TRnC50GrXsJgo8dTGaYIzRlpfSQV7jNfAq/MQkMDwjEqfPZmVQxc/X/VD6hZ
73A8UDIymO/zpsgesEvrF2BhDM6YL0T+UiCdQXwEJspnWd+6svVZhag/C7QK
ljeGplF7kowaQHuKCVgAMkR7RnUnvEEQjGqf1ptoLoPMFhMPONzofVjRyU0H
LL2SJq2JKdioq85e1Yt9R3/DOYYwLfc6x0wsgA6jIou6pw7wVoZ3deZzrSt4
jmMx/XPyUxhOKDGetgTa8jVCUnXgeMVolCQLAbYi9b6keG4DhzIAC5t6O36B
kU5XAS+/ZhvO/SJ5/tcTzxAawFUaJ3fh0wY/ky84eXOJ/ELZxN7TyDZM0K0J
z1u/gCAfMnOYPWD2Mw7tAR+IkH+mInAjg1kZABRnwCxoKo+FlEIzBL5620ZP
92dQIOdVs0VIewg1/53Px68OFR9dCcBr49DwwfyvU1C7LVg6FGR3niVu380Y
aa0L6q4/ctL2UuYOZYiIRdXH/mJeit653X9a0CuMooQlgf6oEC8hFkDpzcpi
lQoLHNumRQ2VEZjQMMW6jbXmqRj64PNoVvZTrRzoiGTZ4JzipKFQ2oQf6v2U
MnUHFdiWMv7kNEho+I8bIh+mC8b/MjoA8iUicQeo4VC1+VPiZFjlP3HpAsiP
1/6Fp5aBzWHZ5kOGCMwDLYWamSCXHwScIMmkplNL0+h+LiXuCen/PRpKgU58
kTrD6fObbEbFMcINybfrR3WZmCa+EbhyragAIEWU+35mbBRegj+sZ162dz6i
1ZvcxZpePeBoC0JvgfkgbO9CQytZUas0uOQHJnH3W74RWh7/ZV9Mg5y6g5Yi
YkKqr3YTb7yPqJuK/V4OEzBfdh5eeeMXzc2TuXBx6cD3U/60kELCyhrmRdVn
jKACE6JNRO7LJFRHRbYE2zWONdCAxaSaEktrXEOSR2YdHSr7pIV9xGFc7dzH
aC6Q0k+rQ/8k8Jflw4d97x0+F5GKmEHSpcwNgPPEzbZ2/AeAUirCW0HWJXTd
aqm3cOqa3gNGf7WgtXSVRP6jjz3hoNgDah9MpBKDjz90vR4kC938Hhg139NF
Mwt0bzPSafAlZX+XgvuHnxC1Fmm0M7xV9BEAqrwUCK47FB7EqqOi1yoAJF8b
MGOsR5eggQCc3qQX++gBcTyQN4nnWzj0ucWzUSoIPjbYIpRB7Ks5QjImZlAY
oeJJsEv65dA2kQ3dOwIfPgKY6cLQrzsW5Odr6MAtGzOUs7+p6q7tb00WMKOa
BhzgtMQ1+sj/p0sJMYr7tZ1TIRh2+XORqRAPVqyOR6bzzzgRXuaf6ttYbo98
qX97MYRnkOLy0z3fNewC77mVJ+FPW8qDZOnbdGY+LSyCBVjU0MH5Gi275Dgi
rX3hvU9leMqgUSIXwQk6Jt21VT8Y/EveXrSGrOMcdR+P7h8qVRA0nBU4+SZR
FerCwdQkP+y6tPOwFaWGt0/fFh8TRaurYIm6nsKe9ZH84VQxcXN9MX1YVQsH
6Tj3d+/oOYr+2Xloex0IqTI3cGpkjsdSysk4IkRzw/3p4YblCuSHiAs21XtL
l8wg+w4MxgOMdL5waj+1bbR8ioUBnt9QOI3rKhDy4w4sUEp9gcIK88zxAQqf
6INJKFwGts6cGngB4yIh2qAnbVYegyibetgXIGcg+O7UtOkvK8f6goS7DEye
JNH8bdFBcNcYnb1I4z+eyXl2RXX4CHeQmTzzc4INTlyRui6dg9Jsp4sYiNla
k/Y2hp6lSB/uhlWBPkD2G/hNaBV08ShMeCMzhcu+MIN3z149i928uhiMY6rv
RuzeaNi5phRgr0PAQ0HQz/4sD75kcs698rhMeG2LUlb7k0gPBkbmIaWOGdxE
3XfYdsNEzUaw2W8sC10/fYfqZv1A41jqVv85PGf2fb0y/mLwd+g0aU/6Zu6d
89mfnn4s8SkRfLvBwkYgOsoDkgpooxSV5LhxgdY9whAOOoedD+Y57Wzm0sDL
YSkj6+BFHUEwwm/UzqGhttPb0P+g3fCQ9R9M19+U/QusBRu+fmhMoPnsUmNL
x8eW1uuy3qQNfuVHtdDhsGUyJEPWSN5Bl9mK0qjydcaH6b3R1WMGn/qg0aIT
gxNNFTziXQuZqhUm3pusDjLp3Yh4OlRbj/ed+tfgUIZNfXaAOlyCRGCGk/EZ
AxZNLed3npJI/uBzG4wigutmgf0sr3LRD5ECbS5WeQizEjeNmRm1Q7o44Vmm
QKG7gB9BZUmG8biExooXS7BP6LRS1PXSu3/flaoV++1LFvGwk5mLzls2ZdAF
WVdn8rq1Qh2lrye6Azz4wycQS8h4MeAf0B5W3VxyvQvbKkACAUzdPpKFDF4m
nyGG7iplU1d37ykegDC81Q+ERh4CrJBBb3rpmqmwsw7eYjpFU8nRqs7XKp+K
QXa4ltfkTTGvGlbjR5SH+gdpOSMhK87o+iAefU09b8oR7rGihHR9NL8J2XLi
9B/PsorufvjVLQrG2K5Pn2364C6WgfkP7uLRdUdwK2XKQJToJrJ1iQbzX3fV
yIHqAN8hQwK5iJeawV/BRYSVarIwfzEwTy/nVxGj9S/FNIKbDA/ldPBiycp7
9WyaOpzy5+gLnG6KhfDR+AutjScvSpSDxYY/dZMw4Qjip7qbTHUbnJiq7v9C
UATirfBigWuHBwzpZaV6yOBLY55xffFdJ5/S5qX/F40TfxNsVVM2beY/1YuA
6A79QUpyRUn1QhJDArlafS4RFz7+lrexeOR6U6jB9c4EVmxBfT+7KhIqzSow
7SN85BkhblyF4gouDnLmLb3j5rZRJ3w2pABh+PYcW6ZRO0kUJcINeCABavWj
hQgYm1jmHq4WeLw4qhL2mx2oMNSlwj3dGzui/TUq2zdwMU3u1PVOLOvUEaNv
8jCxsDezRzwlfrbHfWZGocBk+CHmxL+Mcw+X/qt4kDN3/nnmAx5gdcQxpQ5O
fkH2ubZnveqkvyzr1iWGM37MW94iqBz8TeXx8ETrs/c3MJBD5BdQo9qdSZ1q
P/6BpbagLcqaOVCVWyKPgdmkZpp4T0sSS1tYDRwM4BQ3o2iIvF091RcRLIKH
los6d9ma4JqNUtv32J8bMcleQMnOY6EKyySb7ykIsF2qilzF2Grk/QsrGa4U
JP1cJv12Y+b09+vRxOvLn1w1nHc+GtyVOZV0uInBBtmN3IWeuFZgi+KaGWqI
T3YcX+pkojA8zxRK9j9nBYteX4ue3vFhYIvVqef/djdUDU70QiNjcQ+JKf5R
z4Xbb76qECef5EGDNvCONY2NTMMSmZxzXioqmQnC2t0BobhDu9rEmxRXxtl1
VCNOTaWS3BvYzSGGZ3hgbyMYG2CQ8W6ICPp6MNjNdnUllOpm1scOdCfTr/Nq
E84bLCHgayrgEvKugqdED8InCMOHaSS0QfG+hk2ruQEA9wIzY66h3OXo8jjR
8Krzr53zTABzFToW4/rwOIVsopTdQ+s0wOP/bXu4ZpJ2xYCKg89VX6sBHyrT
EEmyOFqUDo/e5BwmGt11cGUV5B8JTQanF8aUaq6I7NmEK0eTcBdrI3Q8am33
Kzd64BfddjaULTNBmrLPGWD/mH5l5Kfh9QFGevwv3M2zC+ct2dizVPEG+qWk
41qO8mnXicBV2EYDJkaSdjgcgE4L2mj86Gkpvhq1sLnnRkGvICr+gsQ8o8sB
vrdqx8C94uUAFwOLMBt7BuU8LuTMbKEnNq4brBg6K08XL4bl6eF41cHdT77l
0bXpp9gFc7pyNZzqLYJkjuFPjnTb4fbu+i7aD9P7SsIegLQUHfzoqqWUlYos
E4BCnuTHD3zkS2uXVsnlSQ+rBvPHq4fs1eKPXq1L13woDSEBkzB5VAVXXO/b
wjqtMkrjLhU05eWCyW5vE43ItQhUVpBIJGDJ0tXQde6Z6C5vJyDVAaiYH+Mx
C38EmdgjOvzHWI40D9R7WJEh8Zpj+Q+55RhTFwSUCCuXO8F0FSrXGApcHA0D
8w6ei2DFkNzJTgXUnkAtF4DinWYpmeZQTFk62jX3sbnFuMF5MD5Vz5IdZ28t
mfJwYpVGvRuRgSFzUoNSzoFptkCalFegoTK05wdYwTdvPTAXyyb89Yr3exOt
Wj5XGDRecGg4PThHap8oZJwFyDWUPgGIZqYjT9BK8FohvRD6Ddakhtu9ybn5
1f51GIgUGAA/vDAohJAV8im/V/B1NPeUi3iCLwf/8ru/WMKHdGoZeXr//2sI
JHO8hNTM6fGgr3jSNaOxRA7bx5S1vrHPwcnuZ+Dg568nSK2gSUhBKvlVf8gc
lzOiPx+IjVVTMChTPLHfJXPfiDy0UA1hgBUWK0xBEHAwLj2ys36FW+aOWEq0
+QPuHZ9voP8XHrqLLgc4qjLy5GFvZCF85om178kgc8ugPMT9LX8C0ft+gsZL
tzN6Uu1RNE0iY9jAyy2L2POjimXodaCehwW6olPWBWmowZZzBsSD9fj/gpjx
cPYkczbNk55kWThu+ALe42jwRu0TD/zjNKTIpLV8nmMsQSjqdor6+wJ3XuSv
5PjzdvcX3SiECeCk1kRPHhZ7honXcEBJQlUF8FKPg4pZq+ZPD5gKxsu1oq4n
q6Vb0FSnTfL2UZnhc3ywmrV1BDv6El2Re1pxDPENb2eHzQGY8O0UMzcZbcng
hv8fUfD1gzKK58JTAvaZXKhk8XQs3nR6cASWfur8jeoJfm17CjXog20cW44g
QV/8WdQzIicwQx0UdLSek9UX+1RaUp/gagmWCZsz80DY6qyBcD0XMRNNFLeY
ZIojOGkjnCGtCEVnZ+uEMhCuTuW65y/Ailm3DtBalr8dvuURUJ3poE6nDnmr
HK9nr5V9997Inw8dFt7mIBCgcu3ebXHCsYjZWK6yT8DQhRN3VtkdEARBwbTe
oc5N2BrfQELHklG+jM5MmYXCy1iDFeu6mFxQeZCDRv88HU1Afg3rHNMs81cH
5tXSNO+a7Xz7JzQQ1cuEfeRsgRAv3t+v6SjWZkOU1FN8TBcB380IBreViXCe
07mF4DfwOnCbpMtdKzebutRVGqcR4mZ8YPMR9vZWBBo/rw8SpFkD22JbXkkk
kh1Ei5SAU2KDkRzsguM1x9F4Rr2bB+nF68i4OKfYWtQAg/kL5TpFMuK1o8lq
8QEJX473YXFzyUmIxXt5mdFJUc8+xgbl/GQBBeLAxCflzGZoZeMEfYliG09m
tuuGYbC0n+nzo0uVbxCE3u8lO5x6RA8emosmIbT51+nEJryGHqSixzz9sxtE
QzZK+Xn0WiAuc/7HPRE8+4e7GxZN3/15QcWQR0fQxzTZpBalXJYWpaMSIEwo
gXtmqv0l1zJbJZdlLmQoVmDC9FfzYmus6AkdSLBwSHb9MrzvgoLA58tW4Fsy
R7vD7LZxd6eJMKaTB/VOG1OrCNwP9W5VX1zlwuweDKUtuGbKuz7CEVW0Uaf9
+3JqTZlT/O75XAH5oaPfrErAiAmbw7Ecj3Kix85rLCwG46lRCXDbW0blxuke
jaKp4HySRc4rsML+0VpXi1lJmT8GtfiFJoGgrjdVdgoxIXZakgDRKGlxX2mt
dds1pgeiqO9VX9VoDQ7TjBnTXtC/Icjae2LFy2dhMiXd8TO+LT2GbSFbBeNQ
QmmcGQLGF2AZ+Z5b72wdAY8eBfAogUL1hTQxiY1510f9+VjrUyNeaPwTxoYH
XzcOxXDtaUEE1kuwYj3aZQaRILci8oqs2AS0WhB7834mKKJSrprwaxNhJfHe
6Y+qBUWEOp1aOVPrjD+useOiobadPQFkcn9yrsTNDB61IKYi4LajIA0QkNBI
6Id9YYEC/cbhRn8OGDZT4JmA82vPqXl19g/ZcZDV7vjRLHEZWzV5r1uPC/gK
+uIhImuJIaSVcTLYYLzSzcX2YsnTM9QrOrhMyGdhRw0nguDH2gEAYu4HYC8A
b+ZLNyOViVrtGf4ApdrVXjPI2Cs7TAP34aPyqy4yNfoSu2DpIamc+vHy01X3
ARFypOxlJUIo7W7p8DNTRB2+14w74bXd9TbpYXzcoQhThW/DJg/bHgjMBJYA
3pMbvplFpsuc3wfDzFSwMEpcT81+GX7RUa7tsrUilI0GZxcoZ47VJolqrm+Z
NgWMecDMTiUZku8QYWrDIG37kHSLorRNbSS056wWw8tkEtMIld9FzB+adUGB
SHP92VVi8/TQNt9lMOtnMyMVvz14RgHrqkpJqecn70hXM2YJo8cMZ7xBy0Fd
hUi6hWyipFC38/QFq8ToM4hfMH45Jk+HEAMP/y7SWUndRCU1fRFxdSFAzCRz
hdQLCmL+syIY+phRgbWT0/kLkCOASN/s0WAFCDrS22APp7gZNI0Jnxh+LIxk
PV0O1yk3rclHS0NdbOpc/l59IY0L0AJFk3V6OuHurlLE2Kkb5Zs1RzHsooFH
ojoSNgRgZpF98KzYLwPLqxxKe47m8un0FBNADGur7rc/lE3w7itq3CtXIb+O
HK/jDehIQmm4l1PQZcVM7EkzxxK8XKcRj3MbGD9lBGUSeEKPm7rCFeu7ImOi
BdOAF7EpOjLhZ8S+6O5VlW3kcSkG/OMsSGgK4xKcjJKqypMkAQPoG0Zsq+IX
NLbm5lPahuV6r8z1JnFBEB2FUPneL0tuAoMUqvSHbav0a9iFCXNS9mJjLGYb
imPF2JCMlTZ6X4rno6ClNbBkNDIhn2lRaY9J1AyWkpe5b/fsh4nGQOF5N5tO
vCFVQvSp+y8d+SSFua2XgxmN9Uvl46tVnv+nt3etVmE3gBoOARe9EDh0q8jD
FjjXJ5Dbvn3/PeMQLehixEY5lySqnTE+ZBOfwRYGKtgVVcSOEvNz0gQFyDPH
Ji4vYJg4hK7swRB3ZvfMslwccMO5OsAT5YVr/kEcJ8sIK+iGJfZQq6JGqS+R
LMZ/ogG2/NScFERHzAEUEM6m900FfcNepD6TD9UdATWqPg3lfWWgnucvPl7F
rJBkhTC12XF5Fa1Bd0hXdFDrXPGWzZnirEteMIN7EjuRiPeKoBXKEO9nxDgh
60n39D9A+oX531sNxNQJXSnkMkeZ84VlyWkVYd/8917qCn9m54Eo9dlJVZzG
pgj2EpEl0raztbB9tAPCtQC4ea0fMnWjFesuGIll36ULxATrrqynjbdFH7O4
DgwHbjfmrXiJ3mksYgCWtc4MKx3jkvHNXWkgWqDXy6swfAX2Itpk59TpvJHn
ZYRBWzjvNWIQA7RB91NK7TnmX16FgbLUALAUfhyFHrIj3aO/Eo52JRKVHc7c
rDBbtkBEISKMBxyZJGIDIlijcK4Zc83juZangYbHVtV9stMUXoARGjCgAhoF
+F7B9TeRFMVRyvc+oozV4ihC/OfigHcQwJZSjqtH1PxbHETfFKZX1NwBr4ZR
A32CCFK3SmzU7ChdgqLc8EyO4a5N+8kknnQ92slnOiqkYekOqjUYExAbq7T0
fzs6+7/WJ4BlVtdVMqElftzwPHMwsrN1o4L01//RYaRFHhouJulAqc8OIuyN
PYa/vvspGUcTCQEsetcv+MVRuhe89i2Lz+cB1i3kOZluRAW/irNqfByoMNYM
PgHCM5iwAWoYI+R5jfEFuSMMSC6DICg59hl3lp3RpB9hsby2PY7qtiv32m5z
2st4Xnr3qIJcstvnWjKZBN/1fVF6WX2XLOyYVCH/LsyEnd9bXR8R4AyXu4kV
TfKJ/ngJa4sLqLbSX8heGUOaiz/zdmECvKFan+yxzGpvwQyjLKJB8dseNeDl
xfADAtp2kkHdd5VdFv25e2wWOMKTX/kO6tAoT2K/vq1eLJxdH24+zJatmBZy
csWrNAWABdsLwjxYjB7HsAAf79scEp6NwNinf6jlqoT7R4Dc5XVNto8Wk5fG
Ky82ALXpLTvK/vn92BNlt/1Vf5XXI4on9brOvutOR+1zGkvocJB0Mhmcw924
4zdY3DLfy5rJttUWKIqJP0e7f7wfBx5nq/KkrPrbG8Ba2ltSOkJu9mz5W1wK
cQHe1czOcmxWoaMQCl76DzrnaoEwMmodSyOF9vdgSxD6Ik269w5krt2VThTr
g+X8wdSQBIdv9UoMlbCkkNLFjbn5zdp5gPI4G8Lov56Pg7WpeG1uyjdATLEg
liShkltNqD3gol8cKONBeNSK2GsBmVrS6fLoMNfW1rHvdCeaoupQemTMquZ/
pLAX/ZBARr5yL174KMw2OJ1ivSvPTePlPfTmggWRY7SXX4wdRGQ2fmWBzzzz
wyXfWKJZUbxcPIem7OFO+B6GhfjqUS2RYhN93Bg8pNF9TrQGAlvIcwahchnm
epQWpawd1qrQzjuQkH0kWWnHOXlNLktcmEyzbiXdlHeCW9jJr2WF4myau2AB
Kwo2cUgyunvzhy5faDEZiKipl66RWxWrArOCKsjJ2jdbArdhn5VcSQf6xpca
SChoxQs8NDx6wn9jNAfHsM0j+DmBSgf0eMDzM+dikI/8CL71yEBtkm2n3kxo
/CC8HLQMYi44oQRKyfH89b+0BpVnGLgwm9T0dVPjS/DnayLgIrlJMjPXbAlB
AYHroGqMuav1rNzKATrB9m6SldOAWgErogJL+1yilMHg2WYZUGHyjVDhqxVc
FCgNonXzwfrEw2ZFr/HmXXd86g/m1RznTC51N3yI/pFC1bqRmsOwHYsY9oNr
vg9tgcFNENeOTOXTPHfd6clVDD/BxgwxmbzyAnL09hVsfzGyVYrvPK91+3Gi
xrepSMVev2widKoyIQ6180tfrWhVk5fW16CLNBtnwup/nK2HAA10QSjCXERD
cFi+FnBM152RKLU9ckzsd9/Nyb2LaJOaCiqs8FIJZbhvfiNu7U7uWj5Nnli+
iF1sNigS263cKE2a9bm2GvncJkRfmDXKu04cTGryxNSCu3g31bxPnPSBOFsC
OgAjPUwk0G2d2gEPK+iVy/vGxdpgOjLqHrcKrsgQkc/IL8p53VjkX+nL0uc5
7+dg5GRw+FGl74oQsSwr+jCrvBMvEfqCcIG4k3LPwc0AX9z4xJA1wjq923LO
7ztxCwFtkRmxnJtAdzZeirjAOTzIQireN4k+y3HYVtbH/KEWivWGnVYOpY9a
DPVzQm23PpPhNDOnXyicrcAjVj59P4CwMvbn3wMkvhag6KxI10fnVdlPqagI
aLbaQnErvc2QgHYNZ+0m84ixK1rKsK9mK8gI7CrNucm+NUuRJV36i7XYM6VB
aFpBH/sZNexd+Ttsy4b50jFvgEcijMsTYXAB0hYxTSMSyxTee7hFrER3hP4i
L4g9WnYTp9Sw2yps7MKB1kHdasmvhGu9cgm4hTinWFFPP2F2QjwLUhMw7gKS
biRr4aBAwgIgeqejZ2ZAZ12DaGkjubb4wqEbWivV1/vOshgCDeJWOUpsmsoV
MMiP+67HLyQYIWnmjXBXZEO1j4vn0gQ8jG/97p+TERL7iUPKYQpVqmQdwP+u
SqJ5KRmP39R7jjoGUed9hEkzGt0DBf5qLY4brsS9KMBUtNN3+Q5HOHPw8PFG
ROGrl7j21JjTkn7USCws5vrTdKfZXGq6DBYZpX5JrYLfPjOOJC3gsMTtnyaJ
squP1qwL/WfP0fznp5VlkWEet/OcyG6sLJyii6VDr0DWSEz/zourqbf5iD+z
Y0Sk7/lqEDuYvrKFsEtvlMjkS+edrMo/yWtyKc5BFU3o3QW31KbngwMKDS4c
ruib4NHtyW2GjgASREDm9M70+pv8tEYadhQlc3mszo6AKVc15jAUyVT9spHU
TcOsWWudjbyB54qD9365YyMWuodcndkcz69c2YCp8H7tDQ+4C3wwxfPerClY
pPP9X0NCHvB6x9z5hBNUxdFepSyu3qRFGis5gKczdHZ8ZM17ELOe8fN+D8/P
c52sOE8IG9rtrSGBSY8uAntMQSUwWLXrwSwJCU8X9UXxboB6YrYVErUOcA1I
utSHNhx7HJJJXtwmbSb+Q30GLaeOTtWQd9P5pkkFHqA1mkrw50GKL/f8VDMm
h1g7ongA/GuRzxwA7aVjh66oZSDDExOw77stv17PFl35UnfxeQT8d+lLc/ic
MtuTR4RXrwfSbbKaj3qqlMJwMOiQHQ/GPHlDFtMKFWcrOTUg3JZzIFOvHe2P
ZZcazT2XJUvVVZoudQsbB/fi9Q2HpYsHRgEXgi6nZ9re4h5D89oC0s0RXqXw
FKFjTfIBq6XslIwwfSKbhM5gALKnewM5ND9cwAfewaUkEYf3erV4Z2ZloRzo
i6wgtxo5hPfk7OnrkreFnCLWTyocL/Ygpngg3Ul1yq/Zt5X5PkJPYoC0GSFX
OMbEvLWuzBEDEwUMBX84e2ANZ9/A3OFg9HZx9oEQmGkCspf1TgZvEZztowSa
A39LZzgXugJQtQI5CN9cz7CikDM93RWJnI4Uvfd0ZH+koNsNDJGSz8q87Mr5
CVTw1q8Se08YoL4bFqR4CRgMgEDULsP4643K+74cygHmmJPzA9YBuJD7HGUq
Bo1qk3RRkywfjvjZ5LShXPtxCFr1VutHwDOdSmkMnibsw0ghpSSix7Zonjyn
dIdbgpShWMvruasmK640DLutpNBFpiQHOgBnL0yDXZdpY3o0lpgo+QZmAIDV
ri0aLpVUOR2/QX6YrhP+XLaaYr6LTJh/JpIH1xodeJwSpaKGaXh9cze8WQWQ
a6txlo03UFPOKBfkai46VjUY8s9N34ZMgEc7fz68dXW39bIiZcX2ZVeXmc9A
ebNJMGK+2bRXTR+qPTkCnEDX4fqcrN012QkMmMtzh3xJa3P3kzoFlQy9YxeE
yApPQVq/XVvw4bWtBznDeKuYULAUF7L+NWzxl4Tv63wIkGVRNvKMeLXLGfBa
RijAL/ti7X4Ch/6A6iG2Pxwmcjy1MqogJP5xeT7UmWvSUfy8ln+ekELRHZOH
m3zSoeKZrTj/R9uMPlQp5pfox+hdJ9DLoHC+mWBxHzx6UrMuvTtW4qbkdOjM
NnAKkXWxf/P/uHIzNadAnjozRokMUO+jTjtjLmVWbjE9OY1DqGgYwIF8Ic+h
JOB8B8SJiTRs3eB4r/Sq+K1QE+X1QcgbuTNCmTm18lZtnrnGDjxjnWIvkYKc
cGQ7kBt1nmynWhGXHPDUl4q0/uOGufLCVd3yWFiNIfFfINZSwhNlqkTeC7aA
tKKFVVoFIcUkFtEz8geWZ76wHXdKRbkdfZp36KOjUAEogTfYrFenWDOy7R0p
+BuIvXXPtYCqxhK3q4TfcuE3j3zDsB2YF5Pl9PdrOgsjtl24qIc/6LgZm+Tz
+DDb+o3S9i/mxG2tmwdizFYJJKkWxpbBwELqspSrwZPWPBnXVj+d1BFNM9di
t2bAgX4HrHE/LNOU4lqmZBsU/ap0ASOQLzvN2SuzNKpfH9BU3uwfOdVzOZJA
K3vUrF6pa+pGIegzaFGJwaHPQPsSDbAoVOysZbgNL1e+FWpxnznraH1veKBG
Z8obvXQQ8kIrpwKMJiG8Ud0xc4RCMiyjQPfAl0UkjMCzyCqfKItmtwymGsLX
0Zzoz2kzbLY61dyy6ack6sbtDAS1ZoGiD4SWFzhLqPCxDkIEjKxYdLskEW2Q
1bySI7BD0LzagelIPJdGDd4VKAy7C6LBTjev6wDRVsssRyLPTcPh5D5bR5Yq
+/NhA0j+7hyEpsJ+wS7Z4fq2SKI3pHu7BfvsM/A7LrJe3m/7ytrPsYAGKdUz
x7TR71eGzpcXgV1vbM9dP19A70BMe0jcE0yz+G6LvzSUdVt3M3GFy/QWwYIH
yLRJKfms608dqDfEE4OscYvmlko0EC1wLhNoUtvFI3PE7i6j9LweG7ooC2YS
EI0M7GF85ec3ihWE0fc956jhBFbFiNsWlwVTESGbcPGqQ1bEpVp2ymnoXanD
AICcjT/Au9ia9qVH/m3kwlU6qRAL3eq23U9BMkomFnEcxtYJL6Nkf8SD89+5
X7tKFtmGanyo6U7ruCwUyhb6nlsp8oLMd0EzgUNkuRdp3PCG2b9GW1VXCCw3
HH/LAbLsUfzSJPNJC++1q7qERctnqKRuGtvRh1e1BtlYStTlRABzYZ94sfBP
ixKFExr/eLhJJf1pAUlO/rOsyBWgkCLXSYMttgLBDsiZoejVCT21tQe7oqWS
XfQqxGUK3NhPFrD/FR1iu7EJaF9dN6tnSxUSYu+e7t1pLSANbm7o7gfxCNAH
gcN64mG7e+sPsYGfyFS0VcmgpmZIbbRogUUImI8aNrKbVxK3D5bHwQGDzOv2
pOjZf3vH76evgzuNZ+wuqxwQsSKxRElzbmUPVdO49pPGJoZ3gRDisH158UyY
2nJe4TvYJADanxv9/45X1vNgMDC6md8HdPoMVpuRgi2Ig2jGYfE/lwt4bSg0
y+NzBbTdBZQUHeuvnO6oJEmRWO388VEiBg2l3copLiPJHU7YYuhAto4kq00Z
SMzUCFopYN1I/TsGAnb+N4hojGLqZzAtq0lf931sMqIVuJB+RVnU87sKBJRO
R2AMF5hlAmEiy+vz+xvIM5PlHX2IiIt1zAvxQ+hnX+YJGmcM9v/cgkpkE60H
Q4r0pFy1HruANZmt8Afg4p2lMf0yhsdpplxGy5f8XA9wzBPEIQP/+MJHJtWs
ae3nh2CErW7l+P2o+9DKVGVbaXSvA+4RbrcPeIt3Jozs2gNR8WcUn+OLpzzt
/jHuXx1wvq0A+nyi2GsEwUaHdKk7U4FJax1ViKsVatMmkoWXw8X8URceNZnJ
DhMFKyNu0au313SmBSp8S8noEUCAjjGbpZSzfOtVc1aj8wOttMumNLyMNk/I
o+hW6D1sWvYkhMlmoeFnDt0FljDZAKfckqCwxJOy5uaPnP4tbN1O+oeje+i2
P/hMjCgG1y2JnSwI+kd46zKkgjchNPTevC94K8rMfPtCJO6aFrmshgfUgd9T
N7W7M5ueLhPkInvRVKEKuriSCZfKs/EI832VKoiXtLj4Yo3okXaYiTpDCbPr
85+oS0oQPc1xr+/IsgrtuEMZEGeJi7Y6nPzi9th0bsycdn/gRujqXeSpLf/r
QU0H6VuE+c9xfXL4VFsDZAXIQpgbvjFoz9NXyhHMAM6xGS2z465MjTfKLmGi
XAzfyhWHfDTuByAqVrf+JxPnk5eczdKHXhbuE9bwu7Q/rOOQ3PTCvwEX9Tic
c6MhNKHg4kUo/U2VgmGpePoPzaz9JvUAzDPoTvLLhJ5urLfrnmtyzr4uBY08
I7feZBnjXX7yVGmtjcfTYObNXsgTiGP/JTqU2K47th+m9I0Eg873igaTvZN3
zRlAR5Z+lvlIbzWdfs0dvqJAW+qvaH0dp3+9jf1WijJGpaqH3x8yimXV1Tz+
iuhFtM/nXmg6VLYt64y8SuPVcRfoV+vMjY3eYYlwkpIezq9/hyEf/YsQtFRK
Of9Zs7pDMhHiihifAGDrw/alzbUq6nhlTsf4Ml6m7b/kJJnMXJMzGZB/k2n4
hB/IAe48w96jJ9oxf5uxgSRGLk3GZmXY7GtqOh/OsrcrPHMnVrcGnF0DTsBc
y3qTPSRHW9pj6KL7B6w81SCDtKHCJ8J9sYL6coalHJcx7JvdTyBA/0MeiQOD
EE8D5ESEB+62wzxGXwHm3k3VeSAinHZokxVObV/uCz/4e2Aqz8a1sHRFffPZ
jjAl0uPo2dtXsBGrMWHvgiQ2aZv9kiYquSEiDY4z5ihnPGlfzM3JoFKoDF2C
7Y2txtaISFizdjkKFVDqccrmJaWk4T2fVQPVrGAMbp7eeRrg3IN3oqtt52ma
NfaFmfBHfp0jUiXdwVKvnxelbZq6/vs+pUbNy2NecUFsm17iabjSSwG9Uf9d
f4Ax6IGaF4zXDeJ1gnOpp8JP9+CndrVaGCimoBxWM+N1G5k2Z1VFfVIGHaXo
IL5VxIxOjyXO/8Sg/BtUuwaM7UVncWQjPXMJXR5xJjAU2S+3cuJLaRGNV/PJ
JJSwQCWvZ3j0rKa0COg+/RDuTP7+R8fSQ88V0O1ws07GV9GQGkCAYUPstI7a
bMwnZwYbg4lHbAjvMVE8YKeRJI/cJssYMcnHHnPRLvoulJX7Yg7YhbWE9Ve5
hmqSfDlima8YcrO5C+r9DYnVp0bbg8pw1uFWfUUX/jrM0UZOD0PpYVm9veMF
mhlya6cVrDigH6yzKCS1C3RrS6JdDWuufKEXNCg9UKtrxhDSORK3ZXwktA/U
6/3Dc3YV0sb4uDCv6pyehQ+anWHeZdKq/8RguMx0lpJ8Atoyyiq7z/RNJx7Y
FkDSBaSl9V4PGouNvbnRKgOeFVv2eJ2CtrpuZ8eQUmZ7TKOWoWNxaJzFIp5N
j/nM/hJ/6qwLZ1OXMJZEo5sBCF0vofb0nYsteFvwJir3j44j1EK3n1P7sWr2
W2D17lyFd1HkN7NF9RMV+1bC2AiZZA71KJXlULvhaSpAPYG6dIJr2GSiH+/K
Gkwyh2g0ZaRqgI2Z5X2Uf2imi+9VvJht2jRKcCCc0FeP62rLYNiS/a7FtSIj
8lfuBubFQXCODdGhaFZkJvyRgvht9XQGfX1pmf1eo24LcbjoHYCa1JeXGNTN
hOMecoiONEqlvTAgqB8+DBta3Ninm0OChTAqWJ1PDWV+S7Hz5N3GBXLaSr3/
dE1+EWx7J46ftj/v6CNPem8DtJDRuknOZlIEtTOkGoHncsbBYK2uYVlLbzXP
nT42qjOjdc3O3W5vfu78vw0TanERisc9oB/a07iS5XYabxXWkyGBPhdDMuHQ
wXXjmhH5Tm+HE8y4/b16lcIwUfBJyFCk5uD/vGN7PmLQW7g32UZhTJMugSQb
7LQWz/8+NiCzKmFMJeA7k5dGqeLfR8PWml2T7HUEABcowNweape3NvgnRznc
TkvHghDm0FCZTk+A3Anu9Pzikks5VUg+e0bvyQFuJ26msSVoCSSccgWzzx0h
yaV+3M43up5YdQsXrrkIg1Yrcl6lk4B3rn7ObCuFuhLJoAZFRNfFYdZRW4he
bjnPpwQuqFlGG8R6CyCzobO5j+UJWfzijK5KTl1Xa/bxghMDXUwdlzLfOvSy
x422sR5NhkjFT7+qV+IqFLU/2HIUdf+Jp2JBbmtwzFGfNf5bD+gObpUhxxOj
2Q+GQIzrOKOa/fUdII3qUg+9JY8j4+jYJOMCd2XXqaPBhGkoc+8l5xE8hVLH
wsFRFJzsN0fCKxjnTD7v8OfUQQgybWxc9b/PpJ2Eqhd8owbkb+ejRed6fH3T
FBObsCjCGKVrL61a6qsyzdnYWyo2TYfc6iLudlgQrB8xjq7AV75tbwXjxrQL
CqNP3QTBAE8pWyIgdtatR6zUHq52/+dhJqgwwdv5HdKNVvV+KTUDo7yJeJU5
GMD7KodKwWQYA9ch9ao39kPNlqf4KV62iLqktbidJdCtT6Xxk8KcIVvk8fEC
mAB5g5FX9Vg/cvVNLHXzTSAYidQirzDoHiZ0c4aqs93WagZ2KKSvw7YBLjDV
PZqjk+NAEXAeliRFYSVWPBax/6cD/XLh0LKmragqkOsxn04LelURfKqe+KcP
xqxXhtSxThTRsKBxF4ggpliSBNBWnjn8AJ4CLjnvIQ4dvDaFQTkcDyLmv6Ev
AhuduBVrWzmK/W3PAtcEmRZwH1m0yypixbRJeKuDg4cLttahRwC+UQ6GxgjA
Gfni+hP5eSmRpBQAvITQl2Rg3cSIBMqbaka5bnACUbS9K/s/qquEfPA0j+8O
Rli4YIHz5pBsc6PE90JtWlNx7eUjic9d0qoqPhl1kd0vkbCApA9OpeO+cHDa
wIkGJTaT7STFtBeeBD/zRvLlkGltbingGF/E3VDZ1++kHL6RdfyVR9U4L32q
6RvWtzuNTdRqxJsg/f6nzHEEJyaoiqvkW+9LRPuLv0Gth+nfXm56Y8ccmA3W
FUmooY5h15J0xfOHYYxOix9m/Fv4fbDhSv0tS8kfkkPVb+N7+B8nECUwmpNn
mC+VUFulx25k+QflBRnh8Ylk4mgTJq+LYoXD14FZeMGea/DxXQelWeti47Me
vauT1kLxnxci8kx1uLHQPvpN6L80vKJ8ClxQjGq8EmftPP5dCfSWfj/BBgWd
Wy9miKR+ACs4fUA2EROB/HAFvz6+e7yc9gdccyV+1BX5rXVFCav9q5FlC9eX
Vg+jfgFZvgB8fFGe0RN9TUfM7QoIG94mTRzpFRUyz4rHVZtool4mP3eMZrPI
c5w1UFA2bNGgj6LuxkcS0MDECYlimZu+iiiaVHzSPmS6rRD4fAKriyIPmjQ+
jqhAY2dl1MBj+Qkx1K+YSX1yUIHC1i7KMNRwdHfVq72/Gsa7xO+e8sj9Yn7W
mXERtZBl1IRQ3tvWCe5Dk3NWiNpYBDo+7U8uti79CndXmhRk1jnYBYwUJ1qq
BlsGSiuij/904fni6aI/4Q5/kaueMoLGkJscwhmONK7Tdhl7KtmZqKx5AbBx
Ux1lW4kmqsmXvDdYDOg8dpc8irOmfF0SGx7w+YblH/kxB9CBnWutB/kVMSfL
f5JlCY+nLZud9W7nAE2XU9pKcFgtPQRr73aHRmLiuJDzmJiv04BCn1o7fGW8
ddAYSmJB+htOJ//oUV8DYvBZ9/8qBbwPMX5r9/AJkG5GAJY4WHboouVG6kZr
QyrMIZ7QvJurNo16Tu6uzJsVg7Ar/qYQ4QadryzODRbhiSeX1IvpLOynGDNm
UwpcGwSCG98z8KBzb+yM4SWKmYp4DZW/SwdLIjqRR8h7O7HDQ65dK0GOfun+
oejYI0tieyLi6CCG6z0QHwn9Hz9aXky3+25C45ydmIoAtqggaal82FtqlYG8
rwhLxUjCtEyQW9ouy3cI6H7FlnfMfgoZPTFYTiOnczYOmwKdEZGTg71N5o41
pKsi71pBJxduvARA0Kp87jPfVCq6dPQMEbOYbQ/Zq1w3KThRr2HatFw0Yaow
LT/NrtDk0Rra3H4Rl4NFZgv2gVSmkTAGbkLv+gucLuQ55DQ9qib423f/7SL+
7H4OYI0GNJwer2yxGDzXZ6McEW2tigPClN8GdSoxI3XFrmDN5yQCzx6I45m6
AJnZYf++wus0GeYbJSHAEreL4rnmygtH/eMNOi29u1lRW3/8tilN2jekPQzH
ilBW42NCQtlYyCggQhDAztuQ/xu3NUsaqIH13H64bAzBqgg9iN3TVYyUM/ip
8phgkF4UyL5GBrHGLA4UCAUcQa3DsO3SiG5GW9mpAr0DGETTC24cMbcevN/z
Wnd0VkXQic2nm9SvJus1cXK03/ld3sn2cc1I6/GerM/Av7AyvR7TAKEBpKx+
KByHEwscLMRf7CnJv4S9hu694QJ42ZDjWj04eNB2XTmq4gHAjsvFP20AZ9aP
i6AUo5UqmRu/epUJLPf7JgwUT3PlhSbu4tDfKB6QPryJNr46ZqzqWRMhQHww
6WGU6r5LQXGaMID0ftVx2zp8zehVdEaUO/XAHokR+DtomoLIZbvp4+Ov94MR
nKjy30ilGIUE/6JkpSH+PF9uy2APaXTor38+umfZyHgnZSHYE63Nix2aB6Dd
DHd25nFHUnd3jAB7TkYgWdFtNcLSknLtzwlKkr5lAUAbejleQBKJ6okWLskw
Z9cqy8IdTaCJTIES3a5rdY8Bjn8940998Vblr0A+2DewREk8MB1Etm082Fbp
xCB/09Ok0a51Ln9wlXYkzwRkqII8Ojx2WDJT0lMvdq4CPCE0su9b7F+Btirz
9r9eMyr2b1OhTvl8jRCQOxGmFltdRaMifweUFOq4jkC3IXOXQDTHljwjDyXa
Hzgwtn9Df6R3XMO6VmIhdZdVFPB+IjCffv+L5bwj+ILCyomisS+mJ5xFOo7a
I45vvq7TF1CMgKnwezAGIInEOFB+4B7YtpgZOabYSmnQuZ8HpUgB15iip1Qp
0M6X+lHR9LAdkIJu5M4HRb7QTh7dgmn6UxunpQzQ+HbIlUhSQAn0BvrMBJbg
+P/OsYQ0FAMq/+Z7xvIjs7lLKGCQFsY78uOcK75xw3GgopI0oFqXiiTbDyFL
ZeXJVwWt4EMQo7F3OtplivSF09TR0F1aUwvInXHIPP5tKNuxIxW45cezFYJO
WTnkMT38ywbuNYJ4ZrzNe92RfSJTGjpgJsna0XMjr1X4G0nq5rs9fBXg5SnC
4uaVpu0F7kjgJPQCuKJx0Vci4hJNP4oYqTyyuAWNbD+dte7g4RG2KI8fzmzb
7ErgwY/QGQGjB1ihQuCZPF9pp47rBkkIx1gr9nmJWYV/Dy+H7Unw1uKIyVov
9Oe+qAVdHzVvX02LleaNDHIvX0c0qwgRYm9iUDhgTxR+3jKTkJxgPwB92YSz
DkNtkdVJQRL3Nl5ZTaFDYvwGlPx4HLU91L1DhI0KnPEqZmd/pTKVwKjkWTuj
nNLJjQac/vSJh+LM/nMqTPd0gSeL2coIuZy/O8fEelB308h0agoQ5uaUmnh/
fGEDzSquFre6aZ3vQNe6SxoLha06mCDfb1D36qOn6Cl/gVY5nv7HkvwRLPvQ
fh0m72WtnqHeiF+GCjSXDXi1vmr6kFvcf6FsoXBwDn1ikYP/7pBjxU3W2XT3
BBWNjO2EJS2pskMx1uqtw7GYyJFeoLbQTg7Y2sIlc4Sy2px/MuoE8sHoG475
wvim8QagnpIfeutVZ7elApD2wTEYg3NCcIPzFwwBAJhOu0kQheY9SFWuQfon
9AeTC6LzWq5z4fuANQ9U974K66yEMlCcPy0lNuBodAG0CunKi7sTKVhyHvkF
32NaE2swY309wSGVnUV2fbBb5nioIebjPdiVHimBNXcHpZmCHNaebaBt3NVI
IEi3TmOmGPx9pfOVie0svsBLhhGaSOrZ8QmXLpGmon77Ig6s7ia4uBr7wLkS
hmxKX6mChb3UPiMix9S3vBet7O6BHsSLnfVNKa7SBYQxDBcWokG/JrHaIjYq
SYGX6R2nNdEnhGiSNg5+O6ZwZHBswIN6a/O3WhkV4fvi+DH0QfJkdtamZc6J
zwdGJhyHYQCOfDIT9aDyNgszgxbADQQWOMjYYO5YBn7Sm4+Y1mHwMdgwvF7Z
2vIqFi7XtBQpf9whX5vYIQQ2zpcMbr1yv8pvnDVkv/bBs8uig0xjX01TNWFI
dDYfFbNK4XwnP+9UoTzD/kf4gfNWqHIXWVqHqqnnC2R+esO9w6RC6mwagc/4
/ASFHT1+lQy4kX0gKZhm8+kcPydhuUoJRss23MjvYu/00f31tTkTvixFLWs4
ah4novp/o4aNRdZOTN74EPZPRJEcIu3n7Y35gk98X5DU6Fidk9OtCRvq3uC0
IfrUcoWJOj0dZcpQoFbJ5mIRzZOB6jVkLXoLq33JitI0f/+rIckvDBSFcw7r
FVcYq0RMFFq5tIWnSQ0EiNgI0IXdejManDVenICdcV4sK5ltM6EFrthb2s6d
X2WtWCoL12nbeVnBecrA4/KccnxH6/he6rJr4aOVOswJmH91MTpW7y1XBR+a
k06X85SmkmsnG0wXlzW/Ix5IB6QsMt88IPMiCoiGk9sJvtQwoNBzOkBJCC6M
gI2VDXVSOclZnO9h68E8v2IXbX8JeXyOkdw284sUbYznE+q0MiQldZj/Aj1I
SXGzenl/rNuVDgOz9NfpoFUVxn0qkO0i0BsAPGNHVfmQH6RS1CWz7aoXTwGE
dAkRsrbrcC/75hxvs48tnqGxBL1qi9K8TG1rKM6UfDPhbM0xMm+S41duuiCg
1k1aCj6ou38ifo1gwyOiuGfXiRm7RaTrhIkK3HHmJdqEJ+z81aGMsbo0VhY9
BDArEqlxP31mV5CHEVsg8OxgdS8p1RyDqbBwSNP3F73m4cA/8Foi9TkeqJ68
H6Hd9kg9/xk/mjrbSO6+8irAEr+LIYZL+iRCtd4GzbE8iVmTm0s3jJTt8s5t
7sLE10/0/d9KOu41tXl8Ix/2yXQLpNNUhqWZkjrurQ2HXTMWNf/17cLgZrtn
5q/ff8SyfDhARBZQUMpcm3t5fAPzuSY9cuDcvE+VZJ8H6evR5jb9GSciqdBK
A64/jZ1hbuqiQeSUjh8Cm7Na0CL6tT6Zfucy+wNLQflKXvnUnqQxOIa9JSZc
6a3v+g5sXGz/KOofhOlV5BH6ReEUfXAKNptApwXkva1ojYPU7eVcQYcV2kU7
C5g3AZj85de5OryRKkSnBxEG+4UuK2WWe8EMfbs1Ns4JsLDJZxrYY1NwE437
Qh/5nXU0K+NQww2mRGaMH9oS94o9j/IuK4PurSBhdNQZS/hEe8GWFuTJla+r
g4aSWqqNluDixXvf3R3tJ9GFEcwf3FUgEfXEbEaB+X93zel7PxXP4HVsl8Em
zX4Bf51/ukmVivyC+aBrwcUSCw4eleUkiA3opJThqj8ZOk54LHj8IwnVJj64
rnQISc7VHqzRXMHg9ILb8rwzHK1RgLCyUJARIs95L406bKnM9l0jj6OTMGg9
N1s0KpzlSJhZXuzg47Rl/E5ojZMBQSko3bj866egf9EVOKmtNX1tbd5FkoBm
gm53rTFYYwGeqRlFT58waNOCP6p4L3XrnScIqCx7pRrklj6lIL56utEpLiZ/
3EWQGaZihAxHbq+N2tk0zWsMbeDiZ5svUTpzyTa/uUwH73rnHjdfDorNoPqy
RajrkIpr8wYQKabdmUsEHwm0krXno+VaV6p0W/JjqrIehGX2+kfYz32ikexk
QFMABAr4q0GfGwvbsyGYcqYF51cYKt2UlXqalWU86nSAIPXlQpAjwkaqS89R
cClgYqyQPJwIbqGwjjbbYqcOZcuOevPpJ6zpQ3f7xUglW343ZDOv/0329zNh
EfAQGeJ9aMFtr4QkAjnA1e5ni0XIMzv5oUK6zuLbFAeT3gYnpGJC2e1IZiH2
STmPiCYjnV/tafwsJW0QsOceeKhAZVio5HieO8wjFSpA7/wx4pG2n32PdnFq
jKi5O9swToNdNLeP93PvEk6QiMvJVSkEwnicsu5QKkhee+DHDeGvVh8awxKp
HV8hZvsRD4+2TbAY5T4V+5CboiNfEoRmlsPmI+HO50jpgsVYvaKfdwX7YLot
+SZgIyF1kAXzY3ma5YNfh+XTaOVJG2B28ab+8DP1k8zA043INjJLlaULaa/7
Va/rsh1i7MwCot3lATmT5HYGvRDq+lokONiDWhLNab08lknRLclCauNyyoBM
mMCyFGuhhgpv7VW8cnTS52XRoYSt0uZ6bp6Wo6KbVBRL9zRuZgBBofnt163C
8R3zIsY4Kpy3tXDAjNX6RGxdMfyIXVnqYrV8UhvNokKS1NHM6zCyGp0VPExy
0P219mDC9rOeF0bTn8IfIfV2nrKQPf25p14tpqvW8O6V7p4BJfp19itTIP5x
b0fJjCVK2NaFKu4TUK4Jzj3/LKwzYVnTCsyQakeg/IsKIODlqrdhlI+3EViv
GNtlYt4jkrO3UsktZ5cqcV48T5nXic0p/eRaJaWqztXUzcD8TwuejWpK9Huh
yTOtLfTBQzcsHUdPGEiST2ic43EVOLLm/713fbVyxw5cJUhuu3tR8VkHSpKR
Ve/NWzIT3VRuvT+57rXHYOcYKfRU2kfW4qt/ZxVzLLTcoQRr61sZ3Gys6k73
bQvVAEB9h6ZPSNcwmP3hvuIVTwYvnK4pRAJGdWWKR1G/y/3YwDAH47sxvMgh
0hEF7MzitlWH107DD4prcdDsAfaW5z1FuatCx+jxH6zHcIrA4g/eVsYw7uGr
GDSRUNLDk3EhLi462yIz6VsX1mGiBMqe6SmecButYhP3lz8+l+N/wjOoalWT
E2iVuLxcHX9DHlaQlZvFu5yzdOeoNPgmtuxwhvBdZEmyUQec1+VRYWxGwTNk
sUq/xr3vdPvCkyYHvxlIRCnCmVPWllvQzMWT++FS/cNnrOQbN67faWxreNfg
MzrHofINJEg7TW6JbvXQIXnw13/h3P4APf0OdCRIinYm2435n38iBjgQTIbQ
dlLdhvS2SnMYkmXblUrNaFFeil4k8lq2Sh+KJdnEgcymoliJncQay8ZL4+Zf
CPUacaVAWt5vqORaB0cAbSfjPSosHu4qw/R2o3THVZ5sgae9Gtyasn4HFtjA
tZH4HCMu6JXQqZ2MBqiJyRG3rHLrTbuCZ/U2SQq2W/4aATIp4Dq4PmTijJei
gZnlB7QVv6pgCs28bN0vEV005bPUyByQEHyKyib0YFzmp1BTH9iONOkszjiO
2xhiFBP0Dm+CfKktZmDbqeEuqLGRmbk7xZoNpPKBHDMRQ5QNz3bXkYrcZSQe
Aooxc/v4+FUqbgau7vXWTowWihqT3VE2HQX4VvIOcvgIlMvryJwSCbgiMlb9
pDXX6QAOL4VxbWWxPwhQbeoz6+Px52kxmO9ckr8z7wJj8mTeJ1qzl8Ype/WT
s3UVeqCAGk6wMsMXQHU5XEYlP5y8oliOPPh26KKTzyZ9RyMmTcur7gstP93I
9KfnNzx80jABKJ71AO9KNcLsLRT6xjLL9hmhCe4QAsnBC+o0rEQWHVHAXVBc
XzhlrerLxSQLuFPny538hEG4khU/WCeeu33/NmMRsd71XraBmuPibhMW8c1X
YjTgylmmYy92DPXAQO/xSzYnRN2zvXUaJF/KWPcozta3l2kcKQp8P6C3lZMv
Krn8Po3RJ+mEflmcA91QGF/3Exea++PxMpECDDs8WQig0JnbSgvl2NIC06fY
OceFDiynviDQEhEui1919fBNE5aVPGctJmSjMldaTdQBn69qnv63rbtzyGLO
2Y4OY6byQFTFmvfSd1GP6Mhw7s/C5MXOPdo/IoMlZ0aYZAubLu9205PpGsVT
FU4AyJBGKAFgsFz4OTV1B2w5GOUV6KyhkIeUf7ArOM+Qol2xaMVUU6+Fs0HC
GTJPH8W+6tYTYn6/mvyvKO8J6xdE9bUX0G0qW0pbIa6M8yEO8EGMoZtTn8VI
Mj1Mk9jQ3knbCyktT0cwi0obubsOVx+aM0+Mnn57K4ihhYG5sEmqd6pdIGpv
iAF/sir4XkTZKM+UHNkjVkoq6hcpH5v/gT/rriGGdU/3xJtdvd254RPmB5++
bHjQBBaihCdzCOH6Mv8laHSkQb62WEfoGe0iSX0EzRzme9OBATEmBJgwbzYL
9JSNkTzL+0AtksPR+seUxefMaKObfvhqshG5477/ixZPoQOjbVrlLlTbnrtH
6NSQRSLNUA+f/uGnN4pNSB8ShgdqSFOxsbSGxo6xYZnEPf94LCGBrN0KXtVm
OSDgG9ARgvDAKhFFGtACEDL6+yrmxpw7FaZdmAS8LGudgArcmf5i0Wb1JSwc
cXhgIJneB9VZb2VOoIO7pZ87vQrZHYiAD/u4UihNLpzEBMfzFa+lzX7qcRvq
skmDeqCpB30spmVVM9gMPZQtwrh0Mag7hZDPN2tVSzkjazoNxaTNC6ExcNiN
43/IDkaCJhJi/AiRMsfY0bXYm91fsAo9OywuHKmNLSZUdkh51HQbwmc9jhQC
ZOVWsWQr91xYfj6Jid1MuQJ0na3Ry0YxN37yzDqh/i7pX2ohJ9rwHwYMD8fq
Qy3eWONyEXGwUyVdmn/qwPpLG7likvhDi1u9JKeP1V1DYKZ79jkHIhcwF4ZB
Ktp5B/hWavBFz96wDf+PNwG6hVdlc2DkrYgWBY81oirAVD+VxblT8twsbCYr
HqDGcFHpeBt18t5qw3jcrc+kzslTGYqbx1EhZYJGG5Z8v3LGkbZt5lq9aC3J
f97YzfJ+LmnJyXBCWXIXWhakb4I51fTAxzL0L6DvZNDledpBiAGORlsx8jfk
ftvXIQjYdCPHfNEyE08hLXNZsJnzczWlSgVkgSHCPGTXeqNaxEJYUqyJwUVF
FasRQ/bRUA/oAsiGSY8WN9sDcj3Bx1TbLVrH0Uea822pd18pJThYumGtCYL2
RCAnJwAm+pIpjdsA3dI5/4GU0moicCPE0J0Jw4kQeB7UZyFc7HAUSuLM/KIF
VSM5407g9n/e2efDqTx8vIBaMKVPLzCjBR7MTk/OoJrw5K12Hn0zCA0fBlEh
6D219I50Gdw7QlYiKi4Wm4kxoBi1esYabBsneWzb6RKeDmHe4jNpwo+7oidA
x4I5GYosMJk4XHWQqrM54SYcK7C1C5DQ89TRS+NMt1RQA6lsNpOXaDFwNcV4
xYpgknE7ftiLy+/dJSUkRGxJWCwgt+k3wSFuuhjtrDeUUGTk02teZSw51t+X
nhp4YzuCtlDM3D6ipVvlPmb4Dfw2Sl5yVNWlMxCystxqgPTzfCkXAgkgKVrM
P3lG9DGTgQ06A+k+QRJR3LJkZ29md5w6f8Tya6bgKUUlg3z6Xi4gFrdysfBT
3vPz7nF9c+Zf4H4OhksDjm+n+TvK3j2TcrGrv+yufv9rGPF8/baZZDrGNeFG
0Rtp3cSPExucg0Sdj+M7O9mRcn0MZOzgJ+WPjZWDIxWCWPJ5/IoGUvS94lX8
aZe6ZsLEDvil+7fYtcnNPp6xxvhRP/foSzyCd2nsMAcThBPLn4CWazzHonr5
Wj3L8U6GUYWboltCYjMLndKKNDBeTWJmBBPAd5hbdXdjMycakr6cHb8isNXb
XZGDdXXLvwOfbyC3GowOkgf7TioSICqMzjoUADRssweMmov7rMNuXqRAaYTG
K6wU4rgWzDEMvNw/y3TMT3YudjNmSB77nPdoK2nWv3tMu4iIijR4i5X/FIOW
YhvX1H+GfvGkrr5P6GEig8HfB2aNmUTOXBfTvqtpPpQjq3RDnWKm1L7RCOWP
yRDhvhJUBqCOEQIN+rylSogfYX5Vx3Yvyxhcur5R9QnQEpvdswKpSzdSLbtP
iFtDRB2ZFf0GJnZ2tEefyqPFb3XNEz5bsFSBun32sD1d0XHS6i6H61Z1PmkZ
mUW6wZwmge9nynxDm5BWz0fFzq7RVt4mX5O7od5KUMX4jB2kPziVE1KlQaxV
a6xu7/twdiIB++WGVOxn1u6nSWihAtBLROVVivWmWTkPCJDz2d6sCqJRgRDf
VFR30Lh9wnveAdiIiHod6ZpbeZDmWDGH3nP/kV6KahM8aO9BdXArGKUAC0OB
3btA2e7OcjfoHEGS7CKiQEFH+jrYQFvUXivIQg3tRXiD8hNMwf+scbAP/6XN
X/6g1GtPd/NcuBZxvthxU4tNTtkfm9g6MUt6ONFpC1GkHm/02NmHqKcGDfYN
/IYMWbI9wuVNJM5KGkGCoxG2xhMhCZKwkHCnybGPanZ7pLfNLExb2NoQ40v2
qQe50B24NQRUS6SKnxSY3JHdiAqIzpTR4Xo2ssJGrqt1+vZZna3/rdageMqH
UQGQ0RFHCpF90Am0oD2lh8qPaMiaKleCzDL7fvePxkHcgreoCaNV/NaLGX9B
lVWqqna6OIcbGHhR8iSjydD93CdoRx+tqVaiiCntBt8ZpnT5rLDDCWG66lfM
osVT3Sgc9NGHl8Jf+zB3q8djnxDNaboauTnyBFbJ4djwoYqSKAU9hpl3TtX7
WaS9ULmHdC7/KjfVjn/f88db4QwPAKYlztQ3G8Rp9S7ViuVfzRxg2P0vXc79
5oonIp9r+RcNA90QGft55gdZ4ichHcEar8dgIqiIaqzNVB0Ri6QvK+iyUg4m
77aARnOTCdEvzbK6L+psRn9QMFzHasisetUP30QoKMTLuUiQGYS9wJzz5jO3
DCNiHPwJPNf7ZD97XZT9Qo9zbT3IQ07YwftqlloVwavPn8kHIqfLYHPvCcLA
uyVWl01HZJrmBpqnaMVghmg27ltmrLnIKnsxLXkXMvJDpcj78as+vuwVgkSL
ARfJWCFV1+ekI5NwsJ3Es8ea3ZBCKn27h77Mh5IGjIOZHJjVn+/neK8Zmkh4
Xx/Ge+PgVPYSuTdUQa/oSpglMESTmrflZYae31hR/3sVSgiy5c1MKTDObeYz
0QrVToyI42GDQmuO4mKHDO4F4JyZKKCU5uRaAL3OIyJpP0WiuH2rMzJNDDGH
iLWuQvi5Azgsx7vfroFozBrKEWCEXwn4WzTV7K84yicsfLKsFLWpEHVde9ZW
FWAJ/BdmEhduaIN7wE+cAMdk3BwMUvp2CedNaixJHWWPoqQwg1WSlOBVGYD3
ugYzzqCJRyTcBoQPuJtOB78JMRSU1jzwsC6p4yTg40GBqRkLn/mauklBfnkw
dk6jVt08zLq4vzbA3bsQR6SVWd73XALD5x8g8zlLG/IwRo9k72HYrhMjuP8F
NF7LGJhk7rZF/psdqOZvXidzIdJRwSSqojEl1fJ3IpBSTFi2hwifc7oUVqjR
zU/e6gu2i5biLmIzDHa8/PFz4vJczsur6uKJqnLXY6op3FWvYJ52yo+BM2+P
Pce2iZ+YKWeBpqxtx+L8MOsRCLY2EDmmA6SxbJdPYF3WseY/GLEmZVOtiUCB
bJ3VhnRiONPIqLrl0MEs/VDeR8DVVklPa18+z8wRkgNSAbaRjP8hL3JHW2Cd
zPcPkEsGusPpYOcJrwPkdPuppntmbA/y/bEQI2nuh5DJhGJWIMdcYeGAD4EC
lNc6F6WFftT3IiLhHXYqjsVOWOkfUhJdYqKjqUsA1ZKnXF5phBuvD5V3iyJA
JBpcNv4N4rLfqerON/EueBAATvI1kIG955SlbgfKAhvyM5LUye6DEU1NBElP
jpGS4AtKF51G5p6SmLMzY9fg2dn4MT9wtFypOwEhvHhffqN4bQkdDqT2vrpZ
+f9LM7g25Bkx9DZotjthJY7JKPUdtDW4h/SmMUKBSWAbb1g52ZUMhROQhun7
x2lBCiZ+FsnuZEJatuEsNLm6t4+zw0em124Is5y7SybpngYfWiEMZjSpGb2J
Om8ofpoxeYoijsOo+bKBwIMqOOkDcX3MPEd082HcC/hxbS3A3oJkH4GE4Khb
dFCZOpFkZwO5LdW3gg8KQDfidPRPSYeA9tk3NG8RPOVFRdQLJEEIKs7SUtnM
kV3BVjsgUseIQLq6BxyhmMFTMfcMIQ+m1siMGBTedlftqmb1RN7WUAp02ZKb
mf55hYZgki9pafdkNle4U3mq6b6EaC+nHNj2F/wfJALqOZpEKQ5x5Sk2+Nhs
ehDbFN5BCJggS2dHKlpWlRsP6BYdsZ2Bi2JndilJ+7bhPsSN8Mhd1hhmGUf+
8TllGRrohP47ufD/V/9qHbTY4+D0n5G/uAPINVNenLQLae0StXCKbgU3lV7K
Unz71mrGAm8eWL6jWeqFm4VvVRGp8Bp1EIEz0HKne77gYH/6BcabrnjNHlm2
w3isGa6OQIEROSTHx3a4b64XFF+RrC5CDYnEP7fElb6YbtHaahIrVoQapa30
p68QxDsPqLiWbniST3BFCul3DDlNp7ERsG92LpbEBdu4PdeIYRRVqX4kH+AE
0u1MTei5IFJIqrJx9Pa2oBhhGAtyEwDGTA8B96JZwIg4VS7J+03xwcJ25+ZY
TptnNO1H00khtjw2+dJbfwScI/fsK6o7/jOcA9v2a6TFcQZIAXWZxb4WuUjr
3noUOSGgSQZY8zeHzyequTScZ58AtOfI7pGcq7FvP3ZxR9uZygX90XC2qLKR
jZ2+dGsF+bq2L7rO0kfHOckAB3iq/UrT6mIoZ4iW/JQzaoaLpiCpS1qES6Ww
Ls5XgED3NHPnCKUpboaUzpK2Okb5rWPL+Eb83IhvcvqDYoSNsZDuXACasrCA
iDkaf7Xkw+DVOJWPCvCF9/a49iKaRUHnc2pub0I2c9SZj+YIPyTvd0sIMIQV
deStNxal8py2uKYMBjXk0L5mGl6reC/Rs13mwSHIDirO+2ZYKaJ8d3O6/g7w
IuOsmp2GPr3fvX2i3qDEycBz5iaeEwMYmjohwAn+pG2CyAO5Bb22oGB0xMBh
Chpo7VKV8Xy/6mrWJSDR8t0iZ4vlN6xNnIkE+YVp9WWKHU1CVyjX1Zo4eJGi
RlXeB7xnTe0pVzT3dukGSqfHhwi1yONeR8K0oETOgU9SRnS1qn2XlBfBr/JX
f8WJnrcG7IcSf2Xqiv14LtM2T8c8Fytfh2eiylrS5rmsj8poZS3RDzp51zwy
3cyrp4UL1u2iShVysIFYy0Cs18oi7clarzwpDTF/wfYUXplYlMYb8v9wKCD+
aBm7kPBNGI9+nqRPUw8RrOjiVHEqUgIS0pc1Dwgnbp90TRSWMPqIVtgEnue6
p92gUdOyv3uYibtXZyHsm2ecATtQaSIloCSRY23/qW1f320XApYD2LXMsBxC
2fEDeCEg4m7HMNvY4vzqPKMFxNsdsUlDz3SmEWk4fh/HagUj4id7wroMxhI2
s1AH6rRptrl2TJ2KgNnG8E3JU83tN7smmRd9oDDvVJNvWejG7Fk6FFSX7yuy
jMIUmf0BEvf8cG9J+imuTHaEeJqRfcTsAHVgdYYPUlpV98eboJQv/SuPT+EE
otxT9YiIuXXQG+z7vqeSkHfVkhcZMJrs0uJoFSHXhQ1lrKZKSMeMs0yTfwca
WY8j684rIPxfziVy7FH1f0vHwdBtYXo1iVAm/KxFBGa/t580if4NxpLZN+QS
1Kt53vihvP5NxjgWqzRo+8jAmAu9U5ezNYc2FYVlqw/bH4YCfeDZ9iPC0AGY
O+53b/JXJciJKlDUTd8a+C7AKQuwLZsheFD9kHpdYZnMSSCHTQfw+cSW4lRn
Ryhfz/NMz2lS7UvAL0B8lRwwfnVal5O0jCdlq3SfgtPThMs87c1VWS3VgNYX
i4hFn4o4OGdpSjT2C4mJhp8oOImPS3FKSMJTy3bvYs1TRgLLUE1mpFmaJe8l
8ul2OpFOiP6lZwKpTsp1YaKCVYnYMm0fYeLLUXKPDpw1qoyyk5fSjd99ZbC1
ssdkpKRwYV2Q7M4D6AAj4HAwGCoa9IefBgd8AQ51WYeu3iG80UTrcoz0X4ph
nMzbb1H334iE+P3g0B0x+1B614Gem39n7VAZQRQhmmw4US+nvMMbK5rDonWf
7DLUFHIv/KEiEV9xtZ9NHprXJB6xzzqiEw/thlrU0R/R5vDKIjxAvolSe+vh
H3nwYH0A+m/lJNu8mvgp1TZzcd80lqZmWuicVbFXMr/btOQXFyDGhlPjzGNR
iG7zC3uYOnJKMahxyma3Ruiw1Tp3SDvN8WwNOmM2fpKEBkQphuEKwc+Qq7am
qCudFisd2dXWHeM7OE5tBas9xDZiEPzuBUUd3Sv6mqcLYecg5hP/KjAttBsx
0s2KAXZkyKOB/2Ze/lW2/BwQe3Lv4PvWA6VD0xm2OJEwfAd64KQ45JktMPMT
LAA2Ac55a+L0Zwmvj1QSYykw/5kH+JJOvJSLLk922w4WXQdWsGmgoWG0pcuA
Wa+hNMcSpZXdfiXuMfq4ik2VeppCUQ0rdAbAO8H+pzcrmCYFLTDUmFHNQZbv
BXU3KlPqFZZGCdCl5ndOUI9HZE3cEgetUan830wm0bWHqK50fOQPNci+Ggwi
EqoCQVQYjbvvOtDJ8dIoHYQhHS3+sakdE8SqgLn4Ff07091a/fE9R48Wpe7G
0y1DrBE3z7h1bhnjxDgUqjjs3T1JG15cfGMW+rqJhqgVcrZNRkbX4kWx5382
V1FKfQ8St4nUw7lB8icKjB78MefwB9fbKL9DWhLWBGZAiWIP9z8O+1E3GsO/
m9OvDUZTWNaDLcc+pdx+lAy8Dz+Wk+Fldt71JNxZx+OsG5BEvwE4rA1jB4W0
8mV8fNd5zqkYOst4MLnrbd3anU+0ejIb3iDv4RrB1ibsXrSigW7kgLRK0Td9
qwVyK2SHbCfAxPmunJ7qVV23ldoL7TZq/pMHNKTwHdOCqPJf5LoSSvRiAL7j
m8Mxkrl7qptN3AMMRCTlz2XWu+vIHnPGLl7k11j3I0pvzqe7r3NCSg2HlG4i
43Lb/aSaMXg4QGmlmCtEy9Zdpw1n01JzAANWIsqI6u9fz1cAbfqfOuh5Yjbd
KiodIKCG/xSWshNbD7JyyDxS3PHOLPZxiTOWduWVK8nGvN1c+92e4s24Krl1
rkoVYNup7E5EsLl2clGlmlYxnix2na4r2qzprETKVo15PKru+sG1Qd+YavWt
Zgbm0Z0UCVKVbjOZPMxaDpuFewmcFGjVM5w0LipqnhMeT7m3rphEEOz9GstJ
1xT2VowSAgo/I15dcH22qDPkS4ATjq88DOMdNBgiX52rQKD9KjPJzVPe9ewG
xlC7C59IhU8eWEUEtikXo4R/zpDFQat+itYOfmrL24AeSOA3844JSDLnZk0I
1+9nzgyEkET/cVdCi78PGT7/T8NSyC3cJ5pvPpZeXLHTGDuKvUyqyl8XPiru
yqyyBFgKZbzf9SK2VTNdvr7TiKw6mwjtBZcYrXfJrMeYcS9hNBsYbnZSiBT6
kk1woQ05U0lMXYrUDhip8e+52oFkHknlEfN9MBlp5U0vxNf9z8sXDqMVMvpy
95OXZtacOJk40iktOdHWqvFbea+eSlXsgOdftfnhvwE+o8uGA6J12j5SAXx4
gIaZRJ366HJz3fVd4eqj7tL4Ov/ctv7y5l664ulkueqoVdx82KqFiKhiOe1j
jo8eylw81yt1fPL4ajRKaDOoKrOT5jWYOSr19u77GpwnZc4xgcEs5LAy5RrJ
oxykN3fzBd8WzQ9/L0N41L4gPVON7yefjfQVkgoQm+cNadeHAOPGaGDE2nPX
duuvqBD85APYaGtVxiMqT+9Ssgwbtvb/66R63YkWZsRcnEgH137d8q8MZRwq
zG7PHlTW/uLPW7YIpm3/8gGPi/sFAPfVYIybLcAW1R5qjAU/GMrsfN0jnSw/
ZCBXCxXLS3uJSmiVZnuUT41GEfKLkmSfgiz3B04iLHRI3WiJHM+JRaxDLBbV
GG1Q+oqtEtyDemgxG1rsWi++ek8ev/5J7Rq7ZF56dz7BnBkxn327JccyinQD
OD2tkQA8WQ2sdDF8UiHgHHLa2thffdBdVn2MpcrZcl/W36zwed2HV6a3gSO3
ZXtNUVoSnvrZKecM6QoGF0129PM82XUAJQWTf60nRJ6rCyCnyRzxhL4t/ogi
U7PiUgi5PdVfw/0pt1e/UjT3LSBydOzjM8XRJ75WWZ26m+Cf7aNWZERcoWM6
pAeENge2WyMFKO6I6KIGPuH666kaTkzj7+Kn3+7QmMUKELQ9Dd2dfn0VEGNM
n5mKMTUWDDkgibi9cKrBXRHQOCkKIuOv0FFysyrheiR1dThgXYJtJ6duylge
F9rmXr/5IoxneM90T41Lx3l3WTZEwYSBGPl0pHtI1dgb32mTvDhbm7EslGVd
3obvXJEZWCe/Ih4QzG13OgwDz+37ykp0u0iDt6czQtEg5gINJIsCvzxkVOJj
U0ZJ/PUnvo5rgjloJ8cuvYquPrSFU0KREJO4tfBv2Fs4jsREW3qGLvrwEffR
2RvnIhjLqOBBWDQi/TuyghpMP0OgbrrQSyCWhvtAvNMC394buqft5Zy98qkf
FNnElhS8KlrRF9DsWzLX1HGOyy5MibLILlAwczGYF6umfENKQApSOfMH3o3x
aBjI7X2NwrJ3iX5v1gkB8AdZMdXAIMmFQ4fYk/Q7t/rr7tSCdRFs2liOIc+r
W0FYFoOzhmIwxXe2OtUG0LRCmVVQ/jE7pxKKO7I3hzPwKnukOVd4BaHXQ9MR
LTynfBi3Ssx5t8EmuEQvFqTb0QXyFva09qxsEh+Nwmp8IOvmswBOxZy2yJxV
/nFrb/rYf4e3rqSQpgj51PiEaXsaSL9wTQMheG48pD7D76aPOJT0ljZ8J7I6
J4hk/DwD7o1Z6KayE4ZPewVaSs4D6f4hvSC66UrEGGFsn10hAOh+R53iVA/q
a4pjGd+hHr1+DOSv1uDgWL6J1qHpB7k6THh0Az/bqcoHqYaO3qW5/RSsUKQk
Ma5p0UvVSib5KqeNmDIVm9aYwOXi8/84jKEcTUx+kNbdzGXdkqtld4ZS03kv
d4j7/1jgThDI0AGVpKK2mfkv3w/EMvCMf7WCsCC6uy7FbovfUJdUln7sD3/E
vpFruuOc3MzGxO8lI22KkyMHFoKGrKgOI0Oww7AB33/4hw3SPpimv7LPQ+4S
eXw1g8Jrh7Lwm5KKFp80mN627+jsPj4l2aZ0Z5GD4XPS0dl0rujI7S1H1yDT
gND4YWcKQ52HXBfbTy1loLpCnQxrj+g3EjBacxcrrtUQJh1ACo+pOpZFR1f5
sBv4TlSbMVUKFuGi7Ze3kMk2lnyfQryEVa3C57l+NmDoXiNy8qHqgvanrvud
7tdPdqc5OkBigIrltqWQPRBH+32NCgLl4jMNFgAdFN88cwiHd5NrbV6t/Yb3
TtFF76Umcl62+R4WFaRsQ+fSM8TKwlKSoi+g+tEM8y8hbVnj9WhCH9k8dB91
84hpEbeZfeSuunELzfiXLWncMIyOuSMPobimYOJJLvjsYDRwrVXnVsiJnvnM
NAhw4G6vAGEYjfbYk7nau/7F/2eMt92CamQewoUWxahD/3IC9JIu9o+a+K8L
VWAVhvx4IwoCsfHmCg+wLq6X4Y/PbVZhkZNvMuL/sUilP2DWLvY0o+ZXf3ZQ
TSqwvv56yyaL/63TfLT/MuE/rW4D335GjIiARVjKyXS6gbrWQGDGSQPDiTar
NyhRROncFdGiAfjN2f4P/sBl6ydKCcgthAIzWXfGMRPJBQ/fBUxAtc4Tkd8N
OMVoxwi7i8X0M0RpcS4p1VbLTZQTIw3Cjar4EOAX9+WhgVXcc7geJbaB416p
eGCOOViFWYsc5pBG5oZeontrCLIXecJSiMONi0gH/zLx1obSocGLnCFmWf9x
G2tkaLpFjYAEHyh85Z70FnD6eVf2gfriHGnjAHRfk+v0+xpTDVq9GxMePY/u
KdXaM2FMSp3WTUEej5slyAvDsG/mUO3o57+ppAQDg5sSmoPl6Lb90mNZvbBw
M1tquCfSVc66kQVvRt/2yPK/i3xe56A7XzMGt1OtMNCj4dBoH3vaSHJIQh1s
NngPUw+9HvaLtijnCcQTPdO9nMDPuhXGm+dGjKUfs7AQYMzFCmgygsc4ubQ+
gwtkgzAyxoKGXOXCYgi5fzyPEwd+saPuVJu8dYSdZrd0IoEkO8C81FD2LpMx
ofVUSN83dpFJIq44K9UX0a8wu0ntd/wpKGx4M9m0l3HGuoKATOhSrvfbbGhz
sH+ay1mlsIa1kDcLxNhVtc+m/nBG4jCHNn4XIjG1s5EAnWVP0qZUs3Gl1KW1
kzl2tfSP81jzhrNlGc8BKrhDAWpVB8z/xo03+iUSfv8Gjy4mxtyNcwObChXA
mWVAnS2vTmePN6BmDlRb4Iby3QykzfEO0BhEhiH9UECCSxW3ujIWUJkjVraM
wXtWD+/uOchw5KVojhed9H3v9PQlW7+McXRkFfiBzkhktmkM+zGUAmZdziLr
3/FNVbRsfkwEhsAYUf6xQLk3rB9VpzrqnUxsYYYTRUEndC1jkCRmzYo+RgtM
87H+/a/cuRPszu0CrFVCin3cKbYOmfvN1GftVAhh+gy/5k4ooLWLbSl4voV5
vZFt+836ytEJYJr+XO0g8je8CQ4j+EgygOEoz+PZkp7pwBzgC6nbycSx7nj9
vp+TiYw6NFeNeANztyyjy5RpakiOexbjuAcCtOkPCnCm1uybzkijjanew8/v
oBde25WYkZKf25v5TgU036QAJXQuh2xEO5VMEGtMzmIfDMvDelDz0LV0Moj3
S9wZbTi5jZP4VOnNZF+ATSo5lJ5Pocl36lR5ziI78JTWK3Bb6XiIqh0Mfy/o
CSgasVWw51InmBsZQhhzwrh3Fx8YL/ZvuDvOcguB4FdA8CayYMcbOWVmX4yp
S9BZRFIvunGYMxdZKg/aga+72Z0WxH8G+5e1Uwuj5JhJRN/v4QgPYMrdU/95
FULsqRc5lhYd+XtEr64ANRIJiagUEMpnjPsE3TnQsvRUlHs4keRQJ+0dvzow
c57jNxOltsYsE/PdXGUykCDwji7T7jS9mjHuOuH60et3YxrHlPV4ilDc74T+
nfPUX3X9f+aA67XpUGwY/q0voQc/r50UaWNR29AOv+a5P6p/SWvOC0WSkYSX
o5RhBoadWlO8+xhnnUI2bmIRMkGJ4PO+t5PYrVgkHnEBmrmrP8lmi0yivAaw
+I31sGtB/JSLlCWpyfuleQTjugREzT8pJ4hIiumVdgUJH3TWfEfTpUeOgjRl
utAT3MvaCLeDosJmERl/IbvMHyAK2YzG+GCPUnDJSj5f0ly0jw64fvgoF3Zh
cWwS7Uut1WcX4lhEZDrJJU9uq3fXP4zShXQT4nKG8NmU2yPxdB0FqKRzV+cZ
VKBCisTnTWSkuvYR7kZYSdYTRf5e90Dj74B/Esmv/7Kcnsnj2R0TYdinGRLx
kwBoeU1Ac3RevXEY1XiKiSsu2L5Lu/Bp2M+Rtx5e3uJfyqHFn2C9kx03AV52
yOd0XueoIaP33n5PGXrueDIBFtdkcG++9X9viNEfbIqUkLsrGrR5psYcXz5c
uzWqyz8HX049VmSxrrzO8LvqyFsBj3diq9j6LvsGAov+wfB8+hBrwmwyFL4d
TjkM35+xRz3xAhoXE9WlaFvPbKhJzhhTv493Qm94TPLuO55IfpSA/GztPahL
cSq55Vgre+WY51sNFdCxeCwqhfnlZQa/yJLawLAyQA5SK4akzny4Lba+gA19
kyeTijLdo39OnrIZXkKd28PrDDXw+q7EEvfytclpIW+9Bz1SZjT8AjXF0qwj
d46f66DUqIfeoAUceYxI3Dh0hoH+OFBfgih4zIz0zRFSR7enL5aWpdllPmhV
230KsD0QGJXQN/XvMVWsxnOTL33gLrvWUU5tFvsepTMNKnjBUUOrVtTsTpRU
8jkJoAaWocyHXYriDiyVs0pIpOE1fkjui7xT7aMmXFAMyaf6FC8ogPC4Ppwo
1lt4hmYz907ZjQK16gqj/6Ud4uOBaHbV+13fjmMgK+6Ptv5jIwk6d0yfrUKn
qNNs675s4t/Fn0dHBI2Nb9IKIaPvhHxCEoKQ0CbiQyuAg9V0+eX8bqVvfeP+
HgPtuRRo8oACBHi8WJVsD6W6VWNp6PqCp4CBns+Ak/5wwKwkWgN+HNJ+pyrD
Ob0XICKd/nsxwIY2VG0lnvb+BMxYgHc3CbJWsh0UeZ5aPc6LHqQL/rNDcjZA
BMm+AZPPRhSLxlYalvnMCekjPDD1o2X6hKjOGdZmaZ3SRrkWTgI5KEn7ec0e
+CYZvKrNGFI4rDXVhOLFRM5+9bn0PHqL5KcVbhg0O6suwiwyiaa8VmNAdSuI
j6h9tLU+T39p7U9ZFBzXX9B+dyE2pgSEZqWTBC4F5CWKctSpVM+GSuWAn7rf
txn2zDjE5JYjLqCEIGN1H7MSXywKc9e+utTL2Jsp2OdDByWHIrftBVyJb79b
eGHoEFsLZQVJXzby+RY69kmWL8FptS/9oG/xC8Qv+gFp/aWZOqBBGq/4vBHo
OmvddUfdgCxMKiTDEjRxbKzoH5a9CCEzza2oOfgDojKD08JCAhi7l6E6fHgN
8N57RJ5DYU5J10JWkBwJBU/yi9xPj2Szq7qLSItGkjRIMUte5orIcZ2j1/id
v80YfgyMgoGraSrknTAJgDL3ODNf1X8DRMjd3vG7wFO6xJHQy0t+8q1Lrhdc
tVkL89jm8nr7h8A7u6kZF1oGJp4/c29lAtfFSMinOOz65Ulptf3SJM9aYPeW
Z/opwUqq5rNr3i9f7mSMwXL4vWsOSI6DDX4WrBrG7cIbBlHynt+HBRUQPfIB
lFcRHmmlM90RQwjlxGLNFLsBwWxQSVHTDzd3b+5XkdlEqs7JhMJVwcT/2qH/
lGWr4WkRBmGS+ti/oCMV8Z9W6qc/TRF0gxGP+r+Fu3pqcL+Lryzsh367CARM
k6nqGb+TFZxo4n4qXUAu14PiEvkK/yB/Hw0orZgc75gEnXpUBcQP5KqX0eZM
joun194h3fd/DTg3Qn2znfTDeRK9koArI5tzjz7K+ehAqWy755mJrTaLIGEK
K9ZJBlL7QE/x3a1aHLJaAcQ6fZ5OFXCC7TXv3NLJPi57ODhVOMxLk6YJ/+jt
KuAQlegq7plnTXbuYEyHlfOAiLaHutWkMQ4/hQVYzbklCEoWIr1CAP0ymgTz
bDmBy+kjADAIFZuL3nUP39CH+VOY/52iM5264n5D9bs+MFvhM30olAlzYHIz
WVamm4PEIWJSNkMhGqJPUZJTFzkHwUmQW/RA4id+ZCpqfd/Za0+a7ZfD9JAk
H0iYBfYW+G9NyPtOKQDokPfZMqiCPUmOEVvFBoyMxL4D/DrbNAc2JoXU9VXZ
JVNyfYQxvCRTdtYID4uynJ+3tp6fqaXdzlJj84mkAX0tpDBhmYHv43EWR5/2
bdMnU05bvFT/j9zuW8BDCqWsFsKEpaCsvIJw0gqi4vtYFCxpuRwLGGP1Lr3C
pnFAWOUPfXkfDPoXVpQ9mx977zSQIw0c4LDjEQ1qKam0qjji48pYT0RsaIFv
niLun0kD1jfy9IcGn/Vk+TZeZYAlyGYNFJTvzBk3g2ysG39K2PsQOBjuZRyI
dfwh1nI/LwT/VC4f5PRAHd5C7MkEkIjMnrH5ydNk7C+bUfGQuDSdL44I7qiQ
p9q8Pb0g4VodamV4blYEURSv76dMLtFlLODF6ux9U4WKTbJSviU50nqlHHQR
W4czhQgKNj7/Tkkyjt+9uhN7yn7mFer0nkDYqi05vv1h6bSejcIj6QrNyF23
wyVZPzJTD3b3qko+14bZHpmYx2oRdEYgONAt2YD1Z2QBNEzcHfwOIjqhMCk+
KD/VCZ+VO9Fsd4PJjfV/aa7y8PDF6kypyOKvnDRUBsvotXx8dM9bz3vZqg2D
00XvcmreTibySc4OeQTdLwpkUzy1m6c1dD4CyG3jwMrt6O+AXT4N0coHn11k
cQcB+wpOpD7DF9c7prNKhFloMHqAwYcRfeMTjmU9a5pmMLX4mOuGJwVq6M5Q
BQy6eaXrlA5stTWytL684k4TZ6BX9AmO6/bVCF2a+SVCuFST1DyKn+JtmGxh
fj+YIQmfsCSiLxKOAlLNnijCkwIY9pykCHb7KVOfhC8TJaEs4WhQDgr61nml
FscniROiUYM78WqE0lNLc/a+3hb9iVNR45KDNHVqEcENlw+J7TAH9ZEAqSSW
Op5ENr5XXcXxDScbCQNaCZm6MQGH2UjXSQDaO5mEF8fdIM73MwtGPDl4CxM0
E3veclr6VPaMas3EttKPAuKipvEd4dFdxHHapucjYonpE/DX4wYBl5aWjL9l
IQ+A2mRRoH80rUdQBt/4t1LcjyX6Do3Eu8gA3fpWT6NbbIRsYwvjMfl2hB12
lqd0ZCI5EtxwJkIRHB/gUqVmnCwKofykK7ynGSqN/m76arKHlcOo8QRC/Y4n
y6q1a4X5TFTFm1Nx4iQEaFzLRhcz9gk3S4k0qt9UNsbOywQrJqctyUXZCpWD
a+nnr4+6e92cSCOS37miNibQf3YPH8GXS5pRw1TYAJJ2IbwggnOudb/G1GAk
EXwRIkoMNYOwFMfRXTjgmbwwaxKGTBpQFbkd3oqwnAFr5ofHgEoejduU3Un/
Z6opSk59wktJyQENp7iABQzswqyDb8hQdXALfCZ3EmCBYA6tnl86MoNyMODr
ihRRaHPhBFapRPzK3vSs3ncBxXaoM47EJtSDBlzF32MfIdBpM4bJYhJA6VvV
8k/5S1VFYSdFMWmGsWWXfunk8MNpTNnVzaYK0mhHWII1Rb/QX1fjWkX2L8Zl
4Tp6ZTOVD0pMr9N3t/V7EBW8mMMMh9JAD7ZsS7Tx6na5vb5Es6+WC7udf3AE
2nr6QX4yckAu0TgamwwpLj1HZPOzuLbsaYICyfuDYes8xcfdtYZwlETNibd2
W81dZG2E9/aJOftqx/QfVToeDplhSeFn16TqKLZru32t1px2AoNg3GS2PKmn
xnMjb0vX++CodgkD5SbqkZfcKUcyUx5I5ItuZRmTQqAAZUv+fw1W7EauHPni
tPnqhYKn0MSIajxA8ciSboW2LzV0RM2guoH8bylOgqWOpXlre7WgdO+Uq8Yv
MDiuF3ji6qs8mwNLOR3Iz7tubXmyRONI6MHffSeGc0l1jLuEKCjm7b8IuOmj
x8ujthUCXkfr3kVSfZYeihP3MqG0Q0ASj3HXJjr1E9icDa0UtU+qsKcndoVg
M++XscZTwmHQ6B0PBCkW6iY1AeOtb2aeSQfRJTbjD2SzxdbW8m3a96Oy8Jjg
KfA0242rpScbhkbmOzbCjmtmJGGukmIRC2ui044yFA8tnmvQrpXRQHEzB3TK
xrFeXg9/5eFI13Mzg/Nun3UPJLgGMjuuLEh31LRDODm9fQ3YOwtqoT0CXYq+
u5KxByiWRiAxjW7TPpZDsmxYMQJnJVd4LX/oSOYXP3PJcD1dMN7ToUQE/ZJi
uafm/kyRK3WatrPS8XpoVl0gy1J1Ey3mlGuZmncSEZSdAv0PekjJpAcaPOub
PtAwRksD9JHom6OzQuoi/HwBkBNETuSmm6ek6m7CFas8eE2LrGrrxnMPQsj4
veEH3shoMK1OKX4I/KdYCI+RdXMpQ/Sksgi47dKz9QGUXrREGvapdHwtoZ4l
Y0wxHlNofunM1fHfc+37FMr+ihfPocWUSHrELHsEQM+E/I9AyffbwtYbAD1P
BAwkhbZW2yCy0r1vVSRiQAcNY7RYIquefkpQmswhJdvfxIggcoKe59U0VJiM
aBfTPn30wZdnJzWehJgiCsgg2zd1LX6thzwdRjR6FAe/snHtqknJ6Km6v/u0
bh3KZAOcq5TFCfsrjmcSSn//b1nhTOqhVaNw95T/9KPY2xoVM2JTNyAYik8D
pvKRWhIDBurqODr/IaXpEDIvxY+LK51pq6kY8ozFeCyntva7A51ymFSWDiBr
kMA+/eR0lzGRofMT6z0jUARTaeHR7eJbSlA6wsj0Lj1y//YFbXRBZm01mhZ+
djAD5ONzibOK0Xkcw9zqhp2Pb41B4/+mvuqLyB56AT8ASPXOhmsU5CzmRkWK
+CaXDkVod8BmJhws74/rQEaYgLH4nLlBiSZXHuu7FfufIGSaYm6P0VZoCKqn
GS2wSUCpTFjufafJ200xACvByAhYhS8yt9k0DNAM56IpYCRpWiOsTSI7R4X0
+iSZL7PnyUi5keHobA3FeTG6nvHC4qK8i5azTRB2M0SN54k7pRawSMcNuMSL
8NeMknL7BjXGAaZlPnGHICgsaYs2RONlXI+bAPU1iyVPf1GHUjb9HgXcOibt
rxhznTsO+Y8JzpRLG+cb7Uk3RbwEGFOlq+5puGGKiGsSDUWrMLYCAdycoY8T
+41O5KYr6+neuDlO+VXYEkmrLU1AcImDdkn4Go4LlaR6EO7HbPfFA0ZMk0aB
w1fmt9empeNpJnMw2ytK9P28I1iYVmyvQ16dxMbbRICj3DuU/2zX0AxUgVBw
LG5NS2I8jbC+PpXGfkExsr4sz1OJZNE9RHjbM8uwp2JDpsChKS5X65toDupM
EIyQujRrUX70/5nrxe11h6RO1/gPC5dAiRNTHmE2LpL88ttGOLpezLORBEQo
LO8S/cytDwRVxNXLEaUTFrNWlDYYV6nkbPff8XAAqF3QR1GNt3l3tJqEc9m9
i9CFCJYYaNRO5QKikdiFSCEtsPrnJ1TIB7EQGQwcXjv/zjQJrXb++IADTXcR
HlXZ1W/CWsdnie4ysqpGWBDpHnz28u2Yr/4bGU/fvWZQKBXpipuFvM72v/ZS
GZE7CifDRfz0apMioQkxCRcuuwLfbgaTfw/tWX9rwCG3W7HZL2exW4A3qUxY
Zb09hRT6WAyGqBcRwhptx4lhkIxd2EOT0DMYz+fRNpwsy77d/B800QyldlGW
Qkrho3BUuiDK4IgsMqmutgOhCtnsQxI9xIMlbq0Rwp1jD3hJvVpwqXNpmQ9m
c7b7izUcP9TvSu6OEFoDn8rgWJXq2OHSfNG8x0Uh3vOd/orUgmNwGKxGj0md
IuYDj7xAV14oDLaaqQB1DpHgaGPDBhLVk/rh4JSdh/xgUEIR1wX3Tj/olE1/
LjW48FnRbDbR3z1Db53pbOidhFR1UmRO6CgYQhvY+dBJGvt9P6V+yPVrOnUA
6PUEFYUH4Dsj1BxlYETZBTXd0RxRKwxKxXEWo34BOK+g7VBZUxL5Ryzj+IZk
FMRebVIWU+XEl10kzFPMpjRfGcrPfDV1SzIwTbM/3hgE4DWSfvUyPT9r1IoD
XdhdTUIUR0091jBU05kNvem+yL4N+8zKrKQ6MMkSaKi8ivZyv3o7p3v8+9xr
tC65ALpurO9Oe6B9GrsBxcflPptjN1ZuIAXw4a7+syx2yxASn9PlUZ9l0Nzv
jRYMdOiiYjXnqvvebO4E/jt5uEh+ogXtgvU219lt1s63uYWiaeYx67i03mFt
dzCU4gm2ulM9zhvTkB5pB+RC/sgUwLV9iWHRIBjpm7tBQCkxIVAj14OHCj/r
ZSVzaqk67+GLW/4/ByOEs1pUW5FLCy/fiU+ccXyUVOrs5DEXAmTtMzLqLuR2
Q6uL2jIRZfy/BaP43fym3Z50MZzfQBSrbniF8Op6hJXavU3fNX99sSNrZIgC
6HEx3Jjb5HdySMW0Zu1zPiDkhzj9wcQUVfLug2HrmG9guyA4hhKXQ2MqDNY3
82gh0H3D/caCOlEmRleBvGeMMrDkdggcf+Dl42AppYsLvEEB0qSI+NFNggr0
3mEnJPBS4kLdpkkxoT0BQtdOtueHcwvFn+bLWYSSKuTDaRb088EJnWTWNQFE
uKIv1oyP/5IZUwvhCtIRIJPC0TznpVaHfWKT19taUK9sbDb99VblSdg4EFGb
8WNXqLVO6WQUqtj5v/PuYOw39KerKn+0Ua+ws1NrJxEtYu2b7Nq1XLpzAeqX
nJ+DulFPxVn4R/BoNOuXgHGdbN2sKqpPMW2lnc7PSz68YgDLpSOM7bbtuLHW
HwHeI2tlVLS4JuEddO/BvizK0zP5EgwTHqe9A1XZO4320i0lITdfDy0R8jIe
dXu+0iWyio72Iecn+lkkSlta/tk0XCg9fsyYz0ADoNhLe0rPYlgNNKQY3jYf
eJF2ryujCFe21dMeAeqz2BUPPtk0EiK44guLu52BlZDNRjp4VxLB2TXx9oOb
ArFRaebr28TBXmVpcpGBGivuRQFS9Oji7+7fhqfmtO55iXstPSWl2AwxXiaE
qADZhEhnKqvqc6S211Kr9Ai16AZsGygpnVMbLIrrswZOUFgvF9gcXhIRCcLt
rMdlrRQ7qQ4eJNGUzdumfk84EcN93k90UdQpp+0zjEJ6sAeW4XzHAP5ovAfo
wBJu5GcbO8GZFOR7JmVMGqduLCITkvN+SJgvR2fd1jxXiVNd3rAYcj88dwTD
eiWBazKa2lbDhQtyOUlIhB2H3BW2nEDY/JYentLHVQzfwzj7/0J1TR3Kyaba
0ppGhdnCI6wIYOEzu7DS6sY5o6fdHvn4uyUJ6zNAY25LwC9r3CxFQ/lCmvlj
HNKIU51INkf3OELRaxd9ax93q6JPQwda6LQJR5G8QdjyPM7jrqVM1DUQSbqS
w/vpUykeUK5qSbzU0kNCB0ia2VAbcLECTHbGV1R+ZZthgH/LaSREU8B5IvI/
H4cfwHZv/SiwAsmwp5FL0ySKgsZOwZ5y2zn7sGeXWHDBc6fEhh0A9QnXZM9h
h0fH4xWTt49WbePKbE8jbVT6m0vyd7uLYe2IpmYaqen29byanxfSPiQZoOJK
d74WDvJ9B0JEC6aWAaqYvCs7pq5ZTSXbS0iZOt2WV6rkVoltdV0cEOHqe+tA
8mggpP6LcyrYt8pCvnHnEHNxXdXe0ziisdhwoZrRW+9RcI71UjL7gOGnykIi
uoXWjXErIYRxwg4cDVGju6Vx9XTkXJ3hnZG9q6daeu9qQs73ZGaHTO2Qv9Up
RDdaQyyXe0Xbp9xcA/nBjBpD2hNWU45BxlRxScJIkYogw5jUYRid505YWdwI
GS9hMVmWkrXa57KnKqN8fpmhsGKATBWaU/OGKBT2eX7ijtXpFcZKTNKnmx1x
GvJMZaxM3ZrPZWwuPjvcD6kzvwPlfKxhZmGNIh9YiehpMlyww4xRyNqmyhOg
zUKhe0RyHtyUF5TlGPOyKjuXzxPm+EG/vJ+Y9bx4RG4mxvynmN0R+xJbtTtg
rh2srlxsLiiEZTSeCPft4+dSYx4DQ06DjM4TxCD4LCLkQ4vos7kgmqehh13h
4gSplXdifvRaZd/Hq2Zes1w86jEtBh6/mIjwewns0XARNgA+AQBca8f5SiZC
UTrOHAQcxZ7GzDetiWPYlV7NwQfhzCltlKx/jDF3EYwwfgTh+gWGb1HdZhX5
oeuJq0UsXgNOVAJHJMlSWBWcrDF4ss78WMUal80fmGVz25ULhQ8fUjDfca5r
od00tHKRQN7RwBYM+Z6Bbz/vAQ7zBV6Mg5sy+WIY49PDSy2DjznzJW7NBZ1X
pvLGzprKL6HOhs2vsmeIev3OlOMDsbtVO4C5NPncrZ++s4aDx8JtRXutEglW
QwPQC5d4Hei/F534exyBkgWM4zu0Dq5RSWazEMm5BK7n9sVQEFBAxzBgzkvt
tAacTvbqOecQjLPS/Vo4XWGQcjYMeQPpw6X5rWtX56xgS9IHxSkFJKm6w5T5
+wg+7gzstcvniyw2IJlcw5aAU2ou1k/ymZj5Md1pRSdQn165T+ND+MbJR6iN
ZjCKA1qhcdlhHs4Ugp7P8kt3w+jDmEu7zcYZu1HFkwZZ2JteT3lM99dcS2/r
GPJEh6YlBSrRwOoNQpYv1mJ9mA5wn3TFwK/9gXf7uWCQl6AdA8a1FOwPZYNI
CogXD4f0Wn5rDmVoYwQ88jb9Q/agakuVYZfita76X8Xw7BvnURvZCqrbzfIE
9ukkPCNWOVbg6UN/JzpblEO11jgoSHVJM89mwmQPEJQVRf8VKitbfs2hbf/Q
tXNThvfUbuWEwjtDyjm//NsXwz96U0Qv7Ra3StFU5bxOGSuPgK7JraNhQoow
Nl4hIZP+q69XIEJH53QSXeT6jAtsOWczRxkUpq76gWXfP09d/AZNbiL3i31m
vTl/DBsIP+HqEm9OMomGzTn170PFxpCGwk+lLB+rKyeukPMShG3JDBWWdqTx
u8l99I7dhcI14vyKtCQANMNKHSmvU5NriXQwo6J1PJNMHXOdrFuVkgdaaM0i
Yrjeg7U+SvA3HKZlFfsiXvi+LrWe9PsOH30/Lh6ITVsQgAIXz/lR0y79B9PP
9AIr42fxJTCV4ea/TAd9kW4y/kpKf4hjSRJtVJrdFsX3/8mBEtBzYD3kWAL9
Pd0Y6N1/PvXxLUgkQi101mRWUMZKqDrXFlFmi97uCsKPzWWvz+eS/gVAkdtg
py8YX56tx98jUqYnzQThxyWILDOgknz8x4mtL4qI66OZSIAE/+/cgdxvRjZP
zsW9FovhSqT/r7G66Z04IU6XlPgTNARbjYJTjSiD/Kau/hYe+808Xih4Cs9O
vq+EfP8p/zSPlQlFIE+FuXfDz+qNi1sGlD8iz2/4bepaf7SKENbmHp9HOc3/
jirHveviCSVv7SGt+DLXi9GHAa3ezSAz2H3R3stk3nHzHjELQvfpcnMZ3aDX
ypoaDz9neNOLOPBa+jLy+iWpk9/bivQELbS9Rsda55fy3qrgwiNrCJOfDPb1
durN0Se1bsRCTfzMAx7THSTEY1du5scGGmZzxLIGOaelfophQxMuDQv9w0Ko
crNH+2NtFBNZDX/o0IRRMuyCUZQxnOVMyPedCi8wjlDV224Dhoe6FComqDz8
TSqwJk+30VFEme2VYjIWoFDdJTzqo2kAMQ7lCvM7+2VE/EBRDdluFVa8YD0q
d53dHNIytNC7jamLH5UCvZisRhBbxBLOF2MA6tTsfI0OcYJCHAT5Y46hqhdy
oV3nWWjAwv9NLSZkQFqPPaqggNIn3GAG08Y+nmvVDKs48me1HxjplWXGPLuZ
nRtFDuxdkGvleq0/E9XioMRy2rNfSm6aIFg+gb33jl1dbt5s+ESELoeXh4l9
EHRq9I6Qs3+JydSr8guS7vWFTohbiW6JRtCcrNImiVN9dzctCL6lY7J4l77t
ObWclQeOIa1XILkdQww+Who1s6aTO5XN8EKepR4MSmEOiAMgsQliTQ0Qc62/
8dGQWnkqpiXCHeOG/2Rilbc1qcjlFm2UnK5eZ+DFPN1M1CzQFY+f3GAZXNL8
X4SDeTut1Fezhygw/t3X7kbjpC8tXUTpIVaQIxTgwTG1tRwiiUuMRz7ue47g
pwObRxQkNyk5bRTSTkaSMoZtMM6x0m4SrYiWEeHw2tYWNXa6rBLwZilwqDDQ
BaimKfEG9nXq44bVVIOyeYfc3fG5/lP1a+4ReKQ/piI1bs41troILSIRX3Bg
EF13eE3NZqOuomuWLoWES6xot/vFyQ6D/OOBqIDPr1uDI5g4l7jU4fPmlErc
UN78KB3q8KqwOgKBlKSwstGH77tcEHOASgjLQ2KyeC9JDiyCpiW7ZGJQxjK6
TlGAokuNybtTAFrttMxvKB4Bd4BAno/hoWVbE6WkJ6Qblg8Tmnn+gT9b35vd
Gb5ATXHKuth+xhhHMZidZgjbq4frHCjl4et4eXiBI+80mXHpu9h3rx1cd1rp
KCmka6eTU1DRYoDHtp+CqI3nTmTSNy/snmqtD2LOObHfjaAHNr/xdr3dvn/A
SUdYEEiJRWHGNn4VyR913QEfSduknO0cNn+HPa8bE/RLgrFB1hI3d3e8mnT9
pS5nipD0wPdl/PfZ/XVmwL2jxK9xE3ZPUYncwdc6VG/IoJ/9ezr9nr7jB2G4
CL47sKe+emm/wwVd67+hKTsOxW70Ekwijka35I1g+IWKqsy41IbFXy5sm/LZ
1TYurnv21PN0D8G5Hc35wLnGL5ArvH8k0cRGseLrxxhodqjcBaKerPSo4DzF
FQl7r9YJrjk9UrCMvVXShtCsWtJre1UlHJr/kWi4rzlvi7b4sRodFh8Nn3Zs
PHeTwxc5blXMafdlqwhGALkVBKPNEvD1sG+fPUWwkDt3rMPElP6hhvz55WK/
ZZS5A4lR+tzxnAHLufZGcq5aFkVTTJn+BefMyBJU6Mq/U+O9DcKZIMujapnZ
OXLnLkpi+DS2s/nhI4SqyhySbKGzvdEXksas7mmJw79KPYa2Fo3gJKU9wLdv
wr67/s8MRTc6Q9aHOwP1r1RH4sWeqrIHWDHMwU9Ea/lWzGG6SXUGbhzB5Vhx
RJRL7+2tdHElpbOf5+5ZxK43Pguu6auSQznNt92+4QBy3ZOQOIztJCO6YzW4
QQIr7XSZ+NSbBddBrDRG54gp4Xr1Bo0DQqe6+RBPns8Y4NWfDpepo6cxUrMH
Z43r0kNOfw40yeZGN+l0qfMIKHmbjO59l9ad24/OgRuwG8eQ7cYvcnwZwVlt
ArG7RZDXw6b0QJC/d20CSpdvZYepFGDGKGsG9+hnqO07DqwtGuRLPuW8OyYq
+mrD2yz/p2YcIZxBEnpNWP1qCtHcYIadOOGgFYIEnVoI325VmDxQbdsHr1RP
buNbBjKY/1PNjWkklXXPPRAbBkrXFDUFA7ySDRnvV0ljwvxNSaX/sNgYeRvz
sKzIAPE0yNcP4VCL4EMRj59Xa/Vm7eb+OUaVh8mRdVrDaiKKZhgYTh84refL
Eyhvsae4UyXqJ5DjPtHdoKtKLe8aiXigaIlGnqJ58Etu26KPxlQvyyp6+Jgy
lBzcop4U2uiScNvnlshBRUsZPjhFBGxfdbvlmDZYWYCKg0GKwStKb9pod/Cn
cYE6s7QDHkitueiuNpPUD1UAeqW6H+y507XhLuviexnykmrFupqdr3NPGUY1
qv+vttPaFKs2Oqw8kbBimuciqZ8i3EN6jImkB8/wFUjrbbrSWaDbjJ0DEFbP
mOo7zibZaWOl61edimgEW5Wd0szHx6/L1vdDus63JFZmjwAcJN8kc30VvLgL
ecIzGVwQNTMUNxH08hrOodt6eg3zHAJZvmfkPLLiNxSnb61OSY5Ip4Zn7vlQ
muk/R8/U8v3GCfZido2CRPDxAjzLtQFiVtdkPIGPxViPaxwtKtab+DFc9h9w
oFRmMYLgLS5+OiY2TXY7EM0el58/6pRhoQ1nWjfHMzFOTYLttIVmAynwoQNV
3fvwTcv9wt8jTm9ILkFjJi3KthkrYDsaSHFhiAtkEHcWQn5HS0HdCDtqAFYx
FHy1+FJYx5s5zYacK2k1XTuarEm2Qoq1g7oX4RnxZEbuV5A8AFq68RG4XHZp
iL/FxNaT4EUjmBlBsdkb0E+EElYgYCLGCh41RoSfyJ1hrOp/OvKWw+gfvRCT
2ql7070k14CzsuR1+WsEoXcD0Zjw6sC1xFfqncw3V2AG3HzYQwlWf+rgMise
abIqBdjsOEG/eMTp5CeQltsO7JMmE1xJTqZK+b91Jm/KPkOOC5TiNfHXpvY6
z8qR/y53kSv3VplJ2zSDhQLUJ6afXpzbvfRZlXtKGKP4K6lHexjdIXbiPXCI
kY6A4Qpa09nWiqZx1MBka/2RJzQKrC8ShBPQX0ImVtUe7AaHtDsyxy5pE+wF
SRh5bB6ViyaozYntbFULf2gImLdQEyhD1wdm8Zb154E4LWDEzezyvKRaBkZX
30QG8SZG144IHJsxoMM9IOHGRG+COZO1M43SLQm7wQW6EbmV7T/rGqPd8bO8
h8Hr46RDiaAuh7YDK9jUGzqRzvpSay2Dkj6h42JktliSml9D2dixIZkPWEIR
lhH6ASgdaJCOT2tWtJe3/3Dbk1j0hOi7wXyxxutPL214dHa+aM/UA6QDkNG5
7XrdzZWGIwFhC99eaD/adGqQWWNiAbMtyUEfB6jYKsnvXSFQ9crGI9bk5Omv
NKtAHiT9N+pApyctnb0118LU1PtuzCkiYcdvCe+k87sNkfQTXVQorXllR4pa
yU8gCDdRFggfbrOrO6HABwXMmE2Fkt/Xz2RBHwvtMOYF7ZLlGjWny/D9oTMp
4yb3sAGfZyD3j9SKCSpNQQwQj011+u9WAYC5p2l5yHoS5uxIrSwNLr4i4Y4v
0ojRp6sPKVkYin303s7x3QMmtV6pTFaPVDytXvIj7pEM4mp03vxZnqQzlnYx
zzSV3jGtqrHZddSLFURN5qBUlUGzDcGXe1KDsZ/hQj7CKwqqwXcQMpgftyeQ
iWvz5bcJu6kBp3wvWRmgaMTbKWKDlHJNFyYVOt/hcM/YnVoouExM97Gwb198
WhSoSPO2OVBkEbF9uUZqtDckkv+z1BR7IE3t9wqbzlKuCxrMX9sbb3uxXva3
tynosvNBnOFZfOKwGyZG9Z4LMcP0v8zz+lYD6a3Ppo6dbA2vaq/Sruohh0Cg
jyaQmpyFKgH6qRWoWvTxYjbZp6Xu6YVqG10R61wca8hzwoFSjtXbP7aQ3LPQ
Anm4CfyWV36H+WHJ2vOhmkllXvwI3DyqqqzXIUo8kdU+IHN3kScEfE8s/L6u
txc4j5zZoqlAg8ZcNeT9QXU+C3l03n/SdwZZLSAh2MLSRlrwsc1q2uVTJB6M
L3xdij3foLsxAQFma+3FscxdZXnJsu8gALjR+Cuf5GCOqbG8smn1mZdRoXXZ
00SUZDY7PnXjU69kC7zwu48sVqbJl4/TJD4Cl4IBQvauDg0zpsCLBKanI80X
oOaIFRuLWS7plel9dekQcb3yCULxTfUX+u6R8BH82b61HcWARr2eKwa9vwcP
FZfmTbkHDs+otggDW5dJLHX7mRdqZ9N1L1iZZMbVsiA3gX3BBvJnzDcN52/C
u+jx3ycOJnLYcLzyyEib4RS9zSuACrBBcsXJ6bZpGAbGx6S5fvzIIJIk40Zo
cGwpKWzXo7sKFaN72aodxWunM5n42s3qqow472side5pLgJSo3SyTjymClTD
3vM8JxU7BD6IPInVaNyjejofDktjHo5fZsCX0Rthb+708GVjkfpYbkhejxUp
2kX7hm3VbAG0nNLoZ/RU769Uu40GOBCTziKe5c6gAWeHdQJgpsnCIvFaCLLD
B2JQyOZLsrIMK9Da0dI88VqpYaIiCvbDYEemCLFJXOmJz/Wf4DhViGkELzyi
yOZD1qTZC+jBKYdco1DJGNejWqZ3EPYuv6d6wnP5mvxKp8h+PHmN5D9GNyqq
jGUtEl065LR8m2Z0CPt23jvhP2cI0qp725xYCoImRfqgC/Moff3xhCXdl08z
TmrUtGqw4RW93GRSD/RX0J3Kcuti0UZyAzXKj5wP0qV89u8/RYH2ncLVZ01K
oIw+4F8y1M/s+Uqh0tJXA8LfWnUi9E9xhmEbCweARjQ9HVqJhBZvfVJoJJS6
Tj2oyda9IfqREwLFeLa/l2W1u+hUQnCREtpaRIf3h08q9r0MjsY7t373G/O5
iNnlNMLeJJJguew3lPyJbaMlRrVpeqkhA4d0GDhgzGPHH44REHhmKS64UFco
yb9BZ4nHBTrRIUdYAoAtfxQigU1mFKu9mYx+7k8t+c7NeyuP4P4xRhM2HM8Z
IgVOYYkAQ7OpGtjjtwFGGP5BZ+O0Q1oXMAoGeM6W4cEDqNEiIBOslwu7Bbk1
itDIGvm1QjE5Y1u8bCaYgN/Cg5TBQq5zuIH2nT0Xg2OTRS9Y5kc6igPrwl+b
o15nwf7EcdQM5RHZVr7pIxdftW2ftzCmAQDfaMGI6X5dsApC2yC6rYYqnN2i
qDaxpUAkxaIRkRvXEJ6B6iVr8Dwmjzv+Hea6HFEVJivL+Zs2mqmBbZ6kxR1M
FZe/5D0xpIbUyZMZH0esgdwN8+XzBq9I8MTxOKxGX0+xsRYowdczx4VziMie
FMM0B2vM/jwSma7wVmq94nuc8ZQciG+/9THLt6yxjsTttHkKpJccP3+hHC5E
CnkKaGIEaVv6A1zZhPx1zJbRaM1rFaPaWO6VVr2crRX8larXZ3LQnQE0AXoi
3PRSEdjmmKVfJLTtW9SL3PdQDS67/gkcQMVK4BVouhhPHeCfVlVc6Y5aotoI
tv2dMinWrJaPY6PBNkGzvqvCx6c0z8vRaAw18xBgV/w+vLD3bqJrVk2UdcQY
3CIsRkCi47npnQIH6tmjQTRzXq59xbCJiFpy3bgJAx9fEaxjLsvysSAl/VCy
iVKb4soMssNnRfOGagJNM1HcIHSuKlYRoNq+eqyK4ekcsnZhA1pyJc/S+CKF
/xRvcOi3tERWEbelucLNjD7xxz3DNhWJtta/C0ZJgU4OmXjOCZA+zSCc3vvA
PAWyhLww57laPxXAmphIEulEaxd98L0orye0ZwCm52lRMgP50E9dNB7pS6la
y3MnzHyR1NWNxPONJkvlISVlAvyLJR5ytd/CW7hflsh6X0575XInmxbRO0Zq
8je5gfrFxe1G9unW/7aoxickArtIr/TitmqNzgBtLOGli6qfpFhMkV5O/ZgD
T8wrlMGfECMUc7UAsnzdwI2uycZzuukAy78ByL0k6Ryb4tY6YOifXDzsSon/
rsVycwHOsDlXpVIAHwyKoRS/e/FBKtVSzmZ1XGKnNDPL8L9VG3c89FvSYN93
m1pSU2MKoo2ZIzQVGp09tFrAi8nQvC3/aT48ADrKX+ALR/2ojgYMn+jARlGM
QIZf6gII1SfbnW015NidDjmjhOZzPw7mJOoLD2OXq6X2E/ZZhiptQnojnJju
f/dtuOAgbbNh4Kp+5bfDgm/u+WG/VX21NFoVJYGPnndZpuQHSbB2RygBIyVJ
/IriWUy7gRTSzzXQL9WDXAg26GEyC/ip0qxiP9V685n5EW7Csn8twzjzIbRi
LHXEQlSPR2cCroC2dqMN1Fa5OS9Ti9ZLWHoEORcmFxeCBAj7IPRVAb0ZeGD9
wGgg+/bOhWDfo+I21wnNGbwrDvzZ3q+0mRqPN0E03VYeYqaoNlME89sYjiHa
JagDQGc1vaNK+0jjuI3C/Egu8c0vagd0IZONz7Uve4iatnIfhDksRTuDwGSq
/KwCf/ZQJ9C7MII1l4T8etBtnptjD+0s0uax01yiSQGAj1ituzK8YZMx+F+U
QjA5+8sidM2TibX32iWD9ro3ltCqmxCDtXRaV9WmMmk+b4e7+MQdQIkBReAE
n4CtQVqSd/dCEWFgYiwHXuIsHiov+VXH5DH1/4i7pIAAX0Fqotx4zc/9/iQg
W6eAf4b+LrCpL8QOMVoze2vikw9ApemDS0mNXG//7wR2eKjag9AdPHu/lMPd
RMqP4c346T9X2/9G8V+i/IpI8jfTvcPTStsRnLTN9u2GIVDABjo1e/pHyOv5
PMYBeUzAur3E+9D7Oi5b+OgS+3idQK8lisb6c7+YudO2ccIxwU7cux21iBxe
cRWNJSYpESvKZuZV2yJlCgJ7Ug3G08ebXhd4Zvq57UVM9Ymb98MPwrDXR7IZ
If1gpTllkEKwtX9o8GY7HVY1Y2tnErHaUpDWjy9IUDS6K4MH7SHOlrEROVGK
ZsARV8ckil0raSFb5TsbPXQ357ZmLQA0yrLaUJbnEwMm5HJ9C+TKrIcKmF9R
+yA8IMoCfBgwAJG2Db2nhkbBx/kKzokQIxNEbZY0/pNNewOj6XDA0cyUlGTi
so1y0n+pBhyMzJDpLFBqP9mCwBteaXmLdYc/eCAPhR+A1ilzyzAqYCvAeqZT
RJMd19GjJiQ3t3/rdOSFh1FXafBNRG6Nhm4s/uNhC0tq2e+0KGvaK6HgzwMI
DIL8CxzrxEMKIYa5b9qXrad4nqa6r6AhgGPvl6WtPj2rN92QzikoYQ6Or95f
oCb/xuK+hxhJPI9BtJhaw12jBu99edA4aiij3S5MT09Aabi9E2UcX4GjrCN9
sNJSmnzsgF1zOcvvD5fsT0cuGWKjbxTWTwNJQFM14fu/thKeiMhR68HNKjOk
hi990VCJaNnC3CdGmm4own0kCp+r2UensNFwJoDqF0OeG7ObEdhHobzhMnOa
2O1y1vMzUyyXsJnJ98RIRj7s9AKuS5hHJZelJwefF6U+/1OkpEGURZvzyDm9
4bNEsTGC0Vu8VHKiNtXNUdcse8lkwbjCQZm4fH2GMCUQ/2bt5FRe9vs8iDZQ
GsNab4At7fLLylBRZy4kN1RKJlz47uSR6i5uY4BHTtLP69By1rZnVjNI1oyN
9N+kG8ByfsOLcj+7ve/obqHH5esWZmKMpCVUP4gsmANp8klBqSwpuRcfwD/K
3u9AxgUAZmB5eBOZNuHZWwLLZd6AiY7RzpVS1m2nChptX9/Ri15MTLZWus4M
YJeTvE9xkNnn8NrKukSRm45CjAdm7qShsfbVMPknHj8EvMof8yhHSErJ99X9
aAJ/2+yRpMBcy8z+epWc59gGAEQpWUpgfRVQ49alaP8E8dmGW0VbKUav0L7M
GpxMEHzwavWgupHOTF63KE8ce4LFEHv6II7fuLdh8i7lKAQ7bjA88QW2b5dG
KwRhnpUxENlvCg2jlfK4fWij4c7qKeKbd39qtUZM8l41EHm16rOpN68Ax1dS
aOLrjmixAivVhDyNlrWsNtfedwGua7Pa51qWVCFPLtazPmkPnVkJF3LAjINO
8v22WFnf7/DPNlfqonFMEfE5obGNjIRQ4pNBaIr2jVof75+tZkpVhJjXFc0s
qIdhlg8Y17llkhD58BXkxYoKzOPhDXxBXRhR9AlJKJ6KMn2NOdSEDtJgLNY1
vpa57MAafBfmD//t/cR9ANAgufM88PzYlNVDeVsIBUN1H+VCGDb4ozj0fPiM
ynOowZyAKhrArJPmxzZajaDI0Q0yaElqBe0bOlO3mebY9IDwiD5jBFosdrGb
2YzDZKBgoiJSBv8mI8HuuhjsGMyLnL6jTcxwOT/pIrH8nqdI+kM9Hp+9AXEs
3AD1EUP7gz4VAr2vJBAS/RZXbaQC9T/QDfzIMkdKWFSyLxevE7Bvh97iReUf
emefykuoX/VZmLa4DOnXIo+c6U5cb1SNgoeDiZmvPTiMnIUgWMzE4Q4DEnlL
3ddGqimAiz8FHoEZjv7kUYG+2I5gl1yBtnyUCfsmfrwFv42/hx1dOAuyCmcL
+Y5gSezTOI7CoXhms8AtI0WWvZlHVcwiT+B6BbgTHRi5adgrQ567Q9upgO07
5xilrXCzWeJ6jWtFqdE1MN4LludIUD2Mb8hl84gby9qPO6Kn+jdI7SZn20qK
AEZEKXdtSL90g443sFkta2IE7DHL21OY6YOXcM+cvUvFvZWNSasRGhASt67w
t4n+hRYlppixHu42zVwTrLMJ2MrJ5CjvsFTKT7EVbmmy1qt23Zr1lU01utQd
KuYMhLs5elWoSZshvZWV/rlGf1EaUjleS0wuGIUYtxqdOdZjvYdSx+d1xa6j
XxU/p9FCJGmv+GHtypRIo0qI2hc1pdzdobYuYNFHMgHuo9OCRBxkeQiGzreN
aY8pnyhEtH/KwkG0vg8o+xywAza3jjSf4OoqQXGbPrsKmqtiAkMfPWgA/YPd
Ot4h/6EcwdxV53Tyb6bUMQhj5QdatsHhzeBDYSeyKMlQNSDWAGeTpknysdG0
IPFjxrcOVh7tsYbmbDnWgsHhJoes1IJ9XbV2Yqi/wOUCcdDSaRtLdOGxRhp/
ZzquKgn7NrSrrhDuajpwz74GrBAd+ZKZj28iy+pI8K2isMcUtJvsB4e/DTsk
S5fdsoJHw82xX0B5FOcqcEH9zow5a/LyMqniIivXcluCWoIw/NbVB84Gnkqj
XIl7bU2TYFQFwmBUgI39I4LdZp77UGu56L8g/iGHSfE22gqQMIeOLR+DCfTv
2gRrRF0RGEtYzTCNxryVr4wjhe2tdChJSkWbB7eGpe3j2yVsJsk5u+IKbI/m
IQB5uvP0ybCix9/vxUnY9le1i5MYwGDIECG/Lfh8MBWp8qyhc1UTiyL5+djs
w2relGkoCKhl80N49COuT2GtcGcAD7iP1x80PYWnzX0tsilnHYCs0UwClGfk
ihWJVApbGXrmSqMTbziqVGwtXG1vVCfrbfIJRnWdVgHM3ZikObtNUthjmbmz
X/qt41V1OlmnBWanNvrF0zsAnoiC/M/sXvje8LWLILOou807NdICjpFh/DFm
PJHRLzcb02vprsBTPKEkfRR8if3y7aDoK6SVaB7gwigrOiKXO+6Dr2oewNAj
z+4ixOzZdHQx1hEGUSsvOPKbBo/MXOcMgiGtZ5dsG3QSzpK9hT3Hn7HvSoXb
d4fxK7OaceFHPJ/V2Ll2wPNzQJTO5Z7OGd603zm1WSl3cm1Of5K5+sgglsPS
417tDU+AX4Z3AUzumTJ2YFy24Mkm08Jw70EGdeqHTDJSg1/XuaOMwJCpT3mk
EiWXnbAWBm1ghvQ5voDTN1bjJX2iBLp5VJr+1BZjEhz0p12H8PxsefcM7xIz
+qXE29UGF9+xVBkiwQosLRgR/zgiPqH9q2QdvwngxIJFinV+Pxu3Bbg3Bddm
2ovqr2asIu244kPvLRrARbTmGfCBVsOLlXOYML7j3fuYlnTvp8o5a/aMLKkG
nxWLOXpNk972R/NSZWN9nppS5WWdZ17tUliDZ8kBzvw98h2GBPNwoq+c2HLX
x0P3JeLfpRH8SCETV02orugUyQh14Gy6KbuNa0C6HnqUGDltQZfLCcKfkZe3
lYrJu8MP0IuuXxVyjNpyitlplNutdsMNfGcVjia4lYVQFVE+TWVcsX+2feLb
HkaEN1C47adh1nPJc6MKpLp9g3ulpUJvFusB29EMfjzfGflQNSDnuk2sqMHj
BEaHA6D75mGy9TnSA38zCod1zB107FBj41kIyj5IdfsbL01nbkW19v8oVoNu
lvmHMfY2PO3SZNJoFsho8+GfJ64eCVKXDxUYM/vNGxhULkM0mJinRAZTuwQt
G8fsA1pc2dH9OTqrNkoX3skZAfak2c3yI6gtFtQH2ns27ZqI5YJVaSrtt6Bi
sYU6jJe58CHb1HK/TpK0CJiga6G+HtvjJvnT6xikWvGBT8JsekkmTgxIUEOX
yJSbmOzHFLEGaECIcBTOkLR67ZOtMfMis4AiRZVgx3ckYYCfztSKbtcvMjlJ
KtakGLZrDujsQDx/Z/pga2FVhBnIeFzRNnu2HCw8yAuQ9bVOaFd2HvARE1cs
VCh3t4hnzEr+KlfzHESjw290cnZTJvA8DNiFrbGMLzXDJeQfssU7hyhKTKvm
UUAbKFQubJZLI6UawKPvQWEW5D6wbVT21kuJIdmo60QCK7T7SddHrK6jlqTf
6nJ7OoGttBSG6sYml43Q+xQkW6uUQpMKZ4oCq/oBVBqBuRUW5pXYFQH9sRJu
l1Ob5zLgsstfL32J/qyAKEyyHXEEgW45d93EDtywHZrCsLwrUq9peDKFt5Ow
KLt+NpX1Rd2KmhdFLGkg5nR719U4vdUlgNxgArkKCnxrkM6l0dZywej2Qfk4
b8tOxCH/4kMv0QpIS8CA21AMK8RU54O5+xEL2jM4efr72qGYGdwomcARWgmB
0NO0REt+xX8Swl4jMEFWdXVs65zclxjc7OewuIjRPnfLbf9G8KfYetGlYtJH
oRMe4OV9Np+ymsSIaywT3+3HvdXk4X2xYkRahG6Lk+Y0Oo+Hb5IW67osQxnJ
ssa1xSX6Ve5WLt/UGsWdPtxjBlNAfFtQuD9DnQV+bKV3COQPG7TpGaR8BBdv
WvD2fDxt+EFVu7+GlIDcKa8EsldsvA0KxxVNh8vDcaIBUka74kJ5+oHGHnF1
kuZDWEIYA0tQ/OVoPGnS2JC1n2F3cOmYfjA5FMfeNo76rXnr+Afy1P70JPN6
E4htrx9Q9M2mvwdwrQSyO1ZzA82ij0p9UtUBVumh3B/qB1tZDyE9MgiaYZg1
ETMDDy+R8I2Kg1FKv8eQqNS+EYZ0m8IHvyrdAMJBNUhLRi6VbyktjO3PEKPH
0ke2QH/J40zuMn1/2E+xjx5lRDNCy9b/SBF+xd6tU2BEaiJTTgFoNgOqucYn
b0P7NGBMg6kqmVL78YY1DJrw54AbV8zwZBT4HHCT8yoZkph97v+QT/BcxfQj
djuEAFEvjBbYPPPPa1ZZObFh0oBGTv9JF5jdAqpaLb/rF3UUPfI4Bt+mIw+P
9rJKmwdpcPevatiJb1HlB2lf04DX0f+06CggoCLhBQ1GS80NnhUuyQ1vBUIm
cHdwC44Sj19Nex9BVTTPk1ZLBplRsokPKludql9USuZeVWGuUAA1MPQZx67V
J6XayLznBSYAVQJpDcAaBCiL9H0tJsGRcWUhKd97RiCot7166rOOZIRNvUHN
sPjKGvSNnGNeuW244Kfy/Xnu/60+y9PlmblaxxVFrs7nqEqA29GjKgV4FeJn
/N+hHX2QCgv3hwX842fSTk3mq0QUqHLLcELkLf6gUIhPGPB3z5chsqLS4IRZ
sg6NK75pqCCtspDSz7cFUfB7ASXrWF4uBqImMiSw9nBfHJTfJdZ3U7PHgI0J
hTk98SsuqyzBWtyxwrY+omZSZtiY7tA7Hc/gdQ7api+/TMvFA3nTFSLD4FGM
jLORIREnVOYWmmKDkZOnmOZgOP6G8BpAQMVYGcMrVfG9irQiCVZJ3l9lo+PO
qcgS1zxPh9JGqPfoHmiC1mHVDpJn3SCy9j9jU3CHB1PvAGWyt/UnW/+XLyA8
8X8/yJ/CMwf7d3eIyByR77fQaMkFk6EAxHM/baqk7sdYJH9O+e+rQqFtbEKK
iakUy2vmbRTtXuZiXymyt6eumnHT8Pt0yMdvYul241vRvQ61eAdqFyYXM0c1
yArLD2IyNsI2Z+4xaRbrQy9KngWznhbv/LFeJVRUC+HUu0lQctYU4MsxSnUD
L0dhO2RyRCiA///ls8MZNIBFrHRx4VyTzJPrI5HRTXMnDn5RZn1XUzsnoMxl
m/cjiggfO0uft9AhULjqML2yf72HBg0qDob7Hd/SH849KgUNxBTDYxFkxaOo
KrkHd8vx0wiQ1Z7z5JYxbjQJl6rn/j7R0Ebz0ruNUzErCuKxiuYDh2WNykt4
ETpUWnBahDxigCAP8kDM6Bu2rXLg0wH6T6fR5O8K2nOo3Lb9MyS35Mtq7yvy
C+HoUg0W3ThcJHJCCuQ383QHEvhzVefvscMsayBp5f0EWwt1ibaz96oZcbav
pTqfzo0t2c29x9nSWiUoHaUYLcuP0ZgsFzAC8XTdncwwsswEhaJhlKjlYW+b
u/OIr+jEIKp7jMnpcI773canVd6h/3+RcDNeg8DhPJJn96bt8DDvAwN6YSEj
tUcqdbhfF/9sfgZv3pmdt4nkkrG/mGgwIP5/3CNYaEQRrY4loXTbmD3vDKF0
BdR7VxKVrOss4yElEeWQUhcyv9nySbjiIn20Zbi/DGHue7yOHsLIK0hk/0af
icVms7lmyltt8PzQriTcwKQkwlngUEphEnug3Pz95zteOlEY5U4fIqHHayIi
QA57NeQc0DHO2Z1zqgo5dPjhUbV8uyBmt5dckuj+Fzo+QvI6j9wM7xNCMadh
aBWHvB3lLl+7ebz+zXP3aVTOi9xFSK+WUbqUqZWXUlIhiEW5i/I3BDmL5tF9
mtL3MVI5QIT9UtldrLMHdox36hJPbtU8Sck4KBbITMcz9fpTAGUOoZXrvyKy
4l8/NnD85Q2DgW8W4HHrBrKDCbsglVK9yUl0wLERRy9RkUgVU/iJb95Ta+G4
Nl8UY7Gs0hbi27EBM+idebogyp9Kn553AYsEMwBR1usvtg+F0Yws4PquGaZH
OO8Wtj6lxtzXQwpyi+AHrt/72jjDA/bHtkrywLbnH2O9rQO3HXXcVCy1MWxh
VNtItFJ4ycoWOac1e4NnjJY2DpEZxI/zzjryOPD8pY8+qt8czi/qoh1bM4Q1
yWqej0R5P3JL4xvj11FJwRw5g8iDtoEz98lRuzCY4ghPFUcBHyqMmLrA50gV
B/e4LwifIJVf+br/pqnc25TR0xmy5NzLmBavF7ojSYz/nA5OS6VUOea+TfgP
XM7A6DElB/zD9lcw9r83z/v7vPMS7dhKcOog/3zOtpFFB7Z63LeaPavsl3dK
S+5tcRewYAsVrUXOYve+OXeSAXukIe1wjZnRPdMYCkNi1gkR3LZOJw5wOwNe
eWJK0U6lSA0pvnLUTgNkf+X0s0ajbcW4n2nixey8O+rh4gvtE1vKZoy5MYtC
yYhquQiMXcQVKsZ6BSfWd2W5iZyCAijBKIuVqNeBfZahNhlj/n91tZbP8N0h
k4Qg56ybmF8VMhXj3BUvplbSkZM7IXGhh9h2/D3dODfQgO1U4HboCQwU0xX+
ZBq8Eij+YGqEKurH9fc+pWuuGhI4LmOdYl8MMiey29rOa0PF0CEZ7e0WxuAy
m7OdSioMjGrueZ2oOrSqr5aSkZz4LrMvm3s43v13zlSlvVeZisIizSxRkKLx
yGT86j380Dd6YQuIc6o1tnUDYFVWHLE4hEJxOhfudkZGNQpEKbR/Uu8qWFeW
YDYqTe2XV5HGF5NqzNpWfbhdSQ0EQ+yyTq8c3y6OmDO75lkESoWfvchjZX0A
3gDMNHh9vmYscIvyhgCbpCsX2pqDaf0r7hwEiTBXBQtyTJ00yIhrSGcw0wwT
RZ/0TTgFpIVkQOYJ57bjpnmddIULBytsoWL3X4/KrGBp3LVRUpweChID/wvn
sIQSE1MfMfTTVfP4pj7jkvgy2dLgbbRrkCSSMAeqV8s2VFRFnLZrAdOEQeQh
1inXna7HllrxaSWu6+cw0/rmEuC5zp+1G4fnimv3zt8qMVesqom9F9JPy4OI
sBEcK/e7wZsllgFNX4rcLH2wVCfn+AuFMMBz9ZXDrfS7Cw+LQHpu95NtMtfv
1hBNTzpYAR3M8UdB4Fyucq4LZ/e95BjqCGElVOu1oY7M9Vnu9KEks/unRGhW
YlOGT5MC0v+KYKjRtSuoIczR7sGBTjSiLxQyLIEHvqwmIeeRPCuSJ/ujtHmT
NaN0jlNHCzEaX0R86zzPN9vBUj8PneXdRpMyr/LiGwA7VFA+t+woKUsgqFuo
FblGAwOfeZwL9D5vdvoDabedvvrP0LVVSvww0TqQi6rq6Ki4nMhIfdbbJwCX
30hTset5iXHWamfTvvQt93BZo55/ry9NOQx49+6BWjdbxuGheUAsg+xPNaoc
7x+PBkNe/Ju3NAmlIYUlE507rIBrdipF4mhv0/hHOo0NqJiHRHVNOKODIV94
Y2pE7WgKiH+54n71fGBO6skhxml9yDhuVR+TsmwWCYOjVurYdFrUUSs9ml1a
gfdl2AckAnJqmecz8HaiTecTTKtZUYIRhs/uy9JGoOuVC5hIoghi7UeBHtMB
0Ggo/203PRH7dMcjBeZD22sU+s8lWDl36KDBEi5oJMEaEk4d/Ot+ed8QyibX
nD0MCCmpe0zsta5Dfu7YwpVt0CvQ8VM5cyFTzhknnVGQ19KJ/PPruL404u2i
s6+HiW1wtsGaine/pYUzdQd2bjwqeGxOZ2Ty7bwWshhfJ+OcQ2nLhCEROWq7
Snc72dQ/mzBdoqIotiSQNeP9+++Z2+yTOGpKPiIoDbctimc50KLmHdjh23m6
PlbGkH889rteLCa+TfVGGLTvRpV1h/OCzDGl2ZvU4FE9whRygapz+59qo6KD
gM6MqTpZ5i0YYSLDeGlwtCapWlzriDxEiFNlNxy9xbkx8rQ4rux8CiE5bn/7
Y7GHLkjbZviZxqMgqI4mXpmaLk8MWG92tV/wsLuxeusQoip16UeJoEo/aRNG
0awx5AgmSrJJ8UxkEQ3QnP3m5NFlDxSR9Qkk7PhS6GL5XC3fvvXKTg+9jeD2
nvgyqelbdNr8piOupbmXEQkv/ebZtga+4SVB5E/W4fCdUwgwmkSsSbM/E+sn
2zZtDM2kPKb296VT7Ht2zSrZ2VqyqPPypk32cA2AiwplI2bCA8QFn7ier2dX
r3bsWnT+oT8qc96Eda0gn68Hpwt6gcH5icwa34B0EtfaW2ky+FbKTQIQ+iEx
83gDCwtCm7hHfTqFO7pEPdJn0GmR+qeZn5Sh6wfTN6+6KNcE/7NOCHcV+MSe
TnazsUlRUVB4Uiqpb3qNAM2dMCwX/i/7vSU/Zq2sWG19D/DhZkQlYZxaSqDG
qzacBnbeXO5pUDk2F+oP4oT3i8vAGAZ40RCtUp0YLoNhp5UM6IuLyL9NmHrs
5AkYoAPHBamTPwPa74S/ZiQTmnw7aU9VJ85yPtBnlA8V7D5a8zBPEsgwvhwV
EnVinjuAeq/ZywRPOvd98wvkvhkqTeGw88FWtpcF4tlni6bDI7iOn7upZrAi
D8l9iH475pTVF/8TJ3FC8c56I2glBvZ46mNJz6975YKp0rOOBiOjT0pU15Ac
4BbFGqRKfCSM1h3Xwyfw+Izx37+nMD/biX4h9XsgRLiVzGIC+W90+OXZHy7e
qCI5yLdjIXkliMYxTtePtEvN8sBjMXQTGgpatnIuuexoZcaCuh72dGNhh2bB
tN5+tkr7UUKp1lciPVTptfoDAoKg7hiQcv58pGn5e9l2qmcsUTvlCjcD+ooH
a1pPX6vwcqWpGlEox53ymrTHphxgBxnAOkzSSo1Z4bWI0yxTaibVLRRb69Py
GrElU6lkU+CQvK9z0ha8OfugNAghySC6xOFajgTxKieqrnVrcXOny/TRyx82
GYxq3qA+vNfmWyAHTKEfBhDe56xNs/cacoFQWmfl9pvKjmx3pT9bhLoMGVmi
HS2EK0ECZBpsEDCGoCdyOucU3HlsVgd5iXQ2+sh5y3w4h8YpNuf3juINXWDy
6QF0305MNQ3nXzMySUo55ccAEgrY9jefu/p2kRlF8ql1UVcNS+4VNEliQ0Ik
9RxzvCO1mXsK97gzdFTUJx2bSuua3RrVqnr9FRNC4GB9CLDWYe9icj/vBMrO
Nw1H6sOTdSzDpYyQfuBF4FRC3P1kejH/CQKnx0RqUvyme+0THdkOxcM9KXPD
KbXQbzrzhhhISJHhZaU5feVYWf8N5t5nbCSvm+Bws/Glm3C2594C+qotdTyR
eApHFN7T2rgtHNOQ+NP8ITPcj/aA/OC3UcpVy6cbPqV2XuE2WqFzJApZxvYp
5nDwxRi+F6bAPv9xY98nDjPL87KsC74y/cbJPEkNM2/mj6sQfQwLweJsctEw
JAS54Nrsuab7vwB7VbtAiG7u4bZbf6UJ5AuMiDqAHnT9mAXbbnyAwhr/ThHv
qBNJfQU781siX4JCkwNji3s0sZAtV99oUVJ7pGYbo612rY8p3rVO3JOsvTaJ
FumeeqHfhcA/WqJsFtP2qdIl4ASJ9Amh+/qDGMo7B3QpYGenI+QJrw+WXiz3
NcF1RCMRH4XLdFpQSCNzdmObeLgG9Vv1vNEWzNLPb6cUNggT2/1iwbL6yFE/
Um8nCO4Bn/iG8H9nsPtkiZkO7ATdjADeuxvkYpxV2Z4o5yt3luCpHl0Nk5oX
P2P1NcY8Kxkz76+cbN3UdbDMOJ2OnVllzwx487d/gjJH6IznYJ8Ay3L1bym5
b80/jbAaKyaA9FkvXJqyInSQEKuIOBbEUWVJXZzqRqM+ohG2V6UkMbGKVblV
D4kX4uu4oSod/cv+ovirrbYHzFG7mDp9vfXvIpdU0ck6VvNOfDeAcdH6lFvN
GWGMttde7KFGv+G5QwWGEfx/U1kp/LyLdslchQKAnhzYUqzq1+cMaBbYXqbN
K36DIAi/fGNApmteQ5vzPileDSFGlGSxDsF0v/1AYMHKGS7eBNsBk5lbMxCm
qPr5/mgTUF3cThWmssTfpRNE8GP4/R4KKXA174Mg1nk0lXnw/GJ/tVuwUZoj
0c/F8bWtRbOzFLWxZhVQQxRK/lYZdlMaZZyjmb8lrHtOvbl1C27DF/dfx7Q3
nraDu32c+Y/sGCFakxZCzwf1DuOCinHLKEhBhfHssw0YmrdXFJRxI4AlnB6r
aZ25yNwYti3+rUz8T5upgOhIXkKAqKKHbZbdFKt1OwZfNFFAJbkq9vFETAND
GJl2dIDpCGjhpcvaAsNqUJzEZ4cDvMCxwzap6gL7ns1vIuYsklUa3l/Owu2Q
DQJ+cg8c+NDkO8qH3OnJQbeCBy0YYaYVSx3UqkafGjHmhsh+IjJoDj93EI51
H5XkRXUHAYPNXYRKCPpPpyYcstSovzeLUgk08ngNSOZrMLngdEJ9cIgnJIsE
xE2YmZRkACHOr8TBGdTR9Y9RpgcqFC3lvNmolfojkqMskFx4WxnlKp0vcj4X
3hm7RtavLtrSz85Bq0VAMbsdvf/xq+F9QI9ohP7fG+8IMSwzAcmW/Dk1YIT4
LfrFUhcCIbD4TDYqumlQXbOy9GK/p4qLhUNXL9CkoIq77VBRpZ5fdKjwAbpt
87osOQVEz8mQg/n8HIYrJqfpAlMao86w/fS6rNoOYg9Y15NPoRNmdhjYBHTs
7RNqCCzhe+3aKy/EQ5NNaKzOwATL4G6jPctn+NKGQYHvNE3TyeAecihh4w3I
GgEOnTm9XDV98+uGEubrZBdNrFinSMv/OOOMMyJuRsnkrHQQN0pKE7yJgXJk
7HMrTtrq1i/g0x76XhlqPRHSnwCrPf7e7Qo6KBW12Muwc13g+l+wONOS/RAz
g90Vc5QgVcze9yMOyYkQwC/BYVlmaduHbZDgug+AsgZ+8slBNoft9A0YE7Di
ACHkmhzj0PpGY7nW7R8cEb6XyqUdiMJSFtneU3R+7w9JEeJ2wCEa55igIQj8
/4nZadE2q8xLCR6Ka8ch2R+MCmDbRs9VraYjtP8j3geYqfllBbdrPhgA7al7
9UvrfKSQPIyl+R8GcppLr9B+5JQ+1PbwtrkBIFC1ePgdhH0ZYe3QXIqXkF0p
s6n5sLpNHZs113yn179jl4RiB/PKibi8IFQC7MQaAuXQD7rFfO1uMwoU+osW
OGh12iTtqvRLX2JZS1Mo59Y0SVn3A/JEtNzo8V4g9hsihOvPGRfdX1FCCvGZ
1OjvPTRzXes+xbVBmhEOS0AzJeNvGf/UD8hzI3vwo0RNDkooOcCzEYGm/BKB
ZCrf4p0qlYbCif7cOwxaJbliK9hyjx5NiPA9dTCfsp/lEIjfbpcyjpUrUFMa
a209wnIHVzCPzevVkxYHS9NJ8ggKgcWdiBR3sBlcFTEDPkxiurJW6QDaHakE
CCG70I6+C06SuZ9teoQciB5RJyZREhoA2lpO6yvKW5/aVfZK4R1JXlPzh5lS
CbpUzUs9uiWHGmZXF7bW4jW2I5IeIGgkI953mXLyjF9xRRn5d4yW61E+srG0
bMvGzN/YkOJ5ao0FwkEhTEAMhyszJbwqq1bRvWz4OlYu0kkuYH1fwZHvKRMr
LnnKH9kGnFMNKahRR6lY/8Z2dLVTtiTj0CaQRNmRu+b+StvHA2v2UEgRVld4
kcEtdk8kbPCd9bjVBjtfk2HHXgcYmWjA3lPPHpI/O4zczmJ1SSK/QXF4rSLi
b39+fyxz4jlq2B5pCJYHPcxldUIdODECaXbisf6dDeB3Gf+X1AwDiMnx4ngo
JCidC9/vszMKXk2bUGS6exrnfcPh1s/HKtvl8T5op1ImTgamz8lTXN6/0Bvp
U0FQrvjEOCkoqAEYYwTgYjXtMEaxaz3YphLV5UlZTTEktitO4mGa6iho606y
FrOwUgKfg/hDR20KYXlNmkRPGnckCYyAVnj89KpQdGZeNYNx83dClAVRonpe
Tag1v2S8KooKGpn56eqrq5IdTjpT7Zt4sKzL6tsPViV0elIZndno97mn1Ymz
XSQhLbhnBxBFwm4f/Vi9hEMUvVXxEDZuqQyPokk8dgDCKkJqP5EfAqHoHWpv
8SZTZQhNDxBbuRMIdzZkgA+8Mvy3wVwNbY9FYb8230DP7c9Bw/DlzRdBwETG
kZjVsP24beFsvTAQyn0CS2nrPfWmGnnRINyUNDMywrB84CRr4Mf9sDlfqDtr
NBceTs4Volsdgqt/8eRFL+C4lfTs49LPQxEo4i5zG2j9LaHFGXN4WNOox/Gj
qgY6Zey2nQWMehIVtrtHnHrau6dPNJlQRF1L7y2IaP/ULhmyPDvf1p8LoNlz
HUYnL9XOrBtBIBEQ7H0jgdzq9IFKVv/wd32QanR5arne409EA7b+Qqe20Ac5
CWqPdGFbVvL/p2nqGIfIQ30Ep/FG93xEUMLQMxZjO7mZVZ8XKW2i2uCyL+1S
KZQc96Y0FjzFZdmNT8doyxwiWz1SgwJ/rhq3OIbT3QCkwQO9veKurB5lzcG2
xubF5XL7HyhlqX1femmZo5zEXGaNDSJu0+BzDKQkSwrJUtWgyk6K48a89dLB
YWwtJib+oGDxZkUhSJ0MsBjxAlCxnuE4grK2DPhaQm9k4KiVSAzp2RJ0jL9U
HgqZIfB4Mqsh1YPSt/MrLFrlXD0pAAr52awnKqgmQnurktlWgHL5nUgjEvjW
hkhSvARNxeOV0Fde/Q06JK8o0S2hAh96QHLYGP/ZS0xEIZoNPkqchlBBM98y
87WNcONyKxpX6hrtPa4VDPptjN+XUw9LHUkpfAQHrvvQ+gq9WrXz7Ms9+rZ6
nWFfc2n3Hzscb6LCa67boiOwBwmMZRGf5p4+MKF7nkvrTtE1c+lQzEDSABlV
wyzrZj9CTXVjXEXqdfRkIQg5bgnkUtivOHrzhoqTiQswiS/H6arG7Ra9NcCm
Ys4dyGHNLsboRnkY9n7vZxkPMJDLogsGFVSRMKPUpc2VuOt61x9OAKqvesJV
9JBdeqFKVbVfzGYQ7rUWVf245hd0iJKPcmUfsDAGNj1X8FXFZzY14zaLIwmM
SSXAVG/rZPrVJlVCknPhcGZUGuIa3MhjYHISflBKGqzZEut960Njjw/BpcrW
ILz+j4zhxY9cJjlz0K3lPb1cmtpICHwWcXVA29e+sXKfkeO1a5/kmVoRRsDD
Z8BQmm7isENsRcylWluub/WJkQQi7HWW09a8T8gImVUXofAbu6RlD4WfMCXQ
ZzX1qzGl0qEeHX7+yEwqtA4HRfCXsmvePzXDJQxyb0LyYYYMN5vGOqGYnPzB
8/n23DtxItZtRsi8tVUGbpiZ5/vQ5Nt1Ygt2WZNCacGQXOd4RmRnHWoG3fgy
gO4nSPLyahM70HNI1/vOpq0kzEepAf3IW4gByGUx40P0k5rnSRB1h1RdQ1mU
XIGZJx+BHQFvnmmenxm0yR0T9Q6V87rV6JiT8TUYMsp5IHBylKDXxKYDsw0L
Jx+RAxJoy7h589J+cZDa2+OBHtbb88JqoCCRBf0yDx58SJRHoXEOga/Jg6IK
/ikH7Tb6hND4wxIk9kox/5Z8H//vcdt1EV3a1qk+mfV+k9kYTaw1u+RU7lT5
j6CSM3b3Ry7NWJyDX+J4U2pPfUIW4OdqKgeWJU5k8jNx3ufz+uVWc+MHdyHK
R27cyFd6zE6Uop1vDG4uUqXUwttvWtloHMw2ZjOs0gLJqz4VljuP2lAdoTur
RIiQZhEVqvDbzgCPwDWaAOmp2FV047dYJiKmph/wpgzBoa6QZStPALTY8sO+
s9JgS3QOj7qA0S0PqVPWkoKvjSb3OdqsFNMN9DcaYyDFO1nDSDekJEH6XLpV
p9iVnmt7HZUxwRa8zP/ZcZzLYMLRweY6RkUVPf4ODDZ7GwA8LGbcREGuGmc2
g7Q1FuDgf1NI8wSYLVZB8U6erlptA3d8Y9Wh+8TQgSS/yJkIQr5Sht3hvFDO
2AoZEDqCwI/ckraBYv1MKE6fkuvkpKmOCxp+GpzBe8g36q9adMWE3uV4dRkq
mGLdmbXPjIkGr9nGY0Ujnb8dsAYgLMdUzifHxVjjBRFlYCt3zQbwqalUC/Bo
0gmy6PC24BjUINCejCPn9EFblA2U2gKwX4TRC5QOsiyrZ7Bs7GB22OEs2un1
wfA+gd9fc6qHMBF2psTSOMSkhq3QY9TnLWZITPgtJwjSaiZYGnY/oRkrmh0K
1QjzHtY2DoYKszUrdRRzrjHLj5wVMRRtCpig+Px8dGhPlCABFaSBnWo/Y6nr
hqcqT3B4fNvfOreNKjleSuN0Ql+8Sh8MEHqNTTPBWMIP4gQdwqF/C+Ps7ul2
uo9LHVqj5M2YxEHJ0qlpyIz9V+X2Q2Dago7cKIPLPQ8E0nYqD8u89Ru5emt5
L9ui8AxR0dtMaDATF8oUDVWotPIO9uJEAd6AxNPTaCF+7mO/IC7QhAUDgLCp
c22iZNp2RreF4NsfbnQKEp1tXkQdk+64NiRRemk7Nmde/jM8ih0C/mC8Fq3D
4hTaOV6hkMUb9sG6A2XeY0SvFG0r1QYqOnz/xUe6G/oD14Ee3surNoKyCpg2
Vtb+AEG0imyL+KGHUeBXgUX4Ok7NiZ29i/dzSzMIZ5b5MwfYKWDBOsnA+F8z
93tRM2Pfc4lJmBEl9dQa8SPIN+dLzuJZA0prfib8UWMFtUiHq04f7FrsGf+6
HnURgSV21TBhWD8NqHXcyYATqwMbVFNn57x5Uggk2eq82zmhoFBxEqZnFiuh
LLzOb2Daa1+WHE6WXbCSZpev/hs39CTR4NbdrCmhGGmA4viBAlwJZSKojt0N
wUdWqbQhxeMb9pR4IGOMYCzdrxZ5Nf4UIv14B5IsTD1ebn7yrGFwrsi2u9uy
/Ya2z5oJHDN/kwSnZlXeswjS/oYGnfBqQ1RQiF/soZX/Hk8/FS1SAUf2xJSt
VdSeT3NncfXUNZfzol4/XYfK20tE3Ux0rMJhbEtHDxmzGjLrTjsqBTNR6Lqj
Zsu5BSgNSYj/FlEAB40wdjPBj6xzDlIwq/S0g24KzhNc18awa1Hckg8oSc3k
CVcSdqNc1+fz9BdpyYuqLiek8hlYZKMOU0S4eJ4CJchXNSpzDEKBYDsUaLbi
zLP+a4+jO66pCRH4ZTGi9BIPYvzkIjKnge3b4iFMQSi9o8ci25Trl+ZW6Q+r
P2nVDThRUbteQyx9EVo+L+9+Ko8DOMCQa1F0W66ISyQD1N1read0C3xYc4Wf
nnXLSHn0cudErcMSqS6iJrDeR7/FhanRb9trTsOQWT/JaTXvheP+ZOFpmAaI
YNP7/eULWVBNGqXH6G4aCthu9ZdrwMhyh72zGmzNl2T1kxONwDh2OCDwhxmv
3Wzyfj3ISvueYOHo9Oy3ieIcQHb2P5zPqojs2aGHcFIoTMwIkIr8LgPLbG2n
5KPCLyF8okF3Ghu33rPTGPKEgbHjtB2Akk88PSujDqhoK0RADtq1L7L/rT5V
svTkCKFjxPi7hd/TVtkhx/Rxo1jNUKZkpd2BbUF4vVaPS8J4dIGKNFVtdzWZ
MjRUqvH4/e4l2IKXDVSm31IE+AwX0nS9uMTt/kBMe1Ptg0c+bA2BLE8rUnoe
sOOXHbWbs0MA6iDnLKqU2t0IKDKuM4Av6rD0ZIq/SlMftk+SHTVw8ZhhqHMd
fPDAd91pbZGyb4rNJ5Skf2ZtkiDbsJ9PGB6Rmby/qVN+Jk5Y4rl77wKFmAGt
in/D6B2ydErNxgniYIo/VUkMY/XE3TQjQ0wxsaEjf70WHDLPafvZyAPj4jd+
iFUuiK7F8c9DaqkPGGgEPe2V6Kio8Uct2l/4twQHuIwy8SyKKsuae/vCQcD6
yeqqDdxr5HbV6dUuVkc0qQeXevXFHcflWDiLXVdxRHsHHYkxdKEzR2gz08jW
yAfyNkfwXH0Ze+sSJOOAFYoYMPRi9Lo46GmB05dfPkpN9iKfVonGbTXIZSns
VfTP3pGQbl3YYogAUynawDRQW2scRADBYRbFre0c7RQlcPvc5QbojbvCwzmL
qDvHFrAPhQybrECW+g3d9sA9YhRe7v0TZZc2Liav2Cfg8keK2UHRgoK0mTwI
YIfYliz7axXHuG2WstQli4qr7LjyxikWStEys/XSmTQ8QQo0XPfzQrdvoHUI
xRaw5OCTZAQ3u572X/uxQaXGfDxTp85QpXIipgDVQ6WGAnuf1g6EzqxSMs4H
eAjc7vn2t71+nA+x75/+kr5vXIIzR40mhZiKK903ZZpXvhWDmUBTukuL4qil
DIgX4Ifu7BZbdQ0jiTUJLmrD679fvY2FK5nwWgUbWGTcGtO5aXPE94IUKVpn
JqceNkM+Bc7LFElyaY0p2gLtx+tYg1DKTinos3e9s0g7j0IGixs3CkzH1rvE
5quTfzzbUlQhCokOAEVWS2mxt4hhY9NXYy7pRo+T7K/Wb5fjGPHsyJ7Hy7eI
HnExAUMJwCcIxUoQXhSMHcvkA0nE+coq0YCb/WdlpD1FAg4u3/KdGjS3U3eb
+XbHXk6sSNaZ5g2ll6HUMsZXzrKGbft3TRTE9c2jeNozT/cSUWMRhXK495l+
JQOS75lpnkgsI6Fd6cL3/r51O/WTRTzUGgE29tEKj9KFOCHOYcAZ1i7gksRo
VHpRd1aJYryAw6R5euSGe8kBPzolTreX7upZOuTIpQdFoWosfUI/bkMLf6UZ
dvmBE3vlQ2VUYpx/iGs8OAvpXf8zxjEqyISgUwcLb6mTpW6BKjfmb5873hoF
P+bWsiX7XM4dlFCkbKVcnqOzqmhR8JAhTMcXtdbl4FIy7GLK6hXsfxcKiyKu
+BE1E4t5HRoosQj6KbnRpyBRZutiaIVSngXN1DyDx+Ke4p0bVhDlcRhcyq7n
bQXf5rnwplvian4Mncxlk5iVQNJcLbzW9hQFwug2jx1P9qp40MFb/hgIqQbF
ncEhnJEphwaUeFBv370aXrxE+5oOTBYb0Kba/CcQ+0c2P4hpGdpQ6/7MR6SF
Wbda37gq/Ssa4r1vY7lU3Hu7TtMEQms+R3P1XzUipLaSkPBl4K35rl/5L0bj
wugUUkTFLBWZWvlvTVKK9zG/SPs/PdnVqv+xeHdcmWMamc/S5mpNgnBVdVXS
SXPmrog/7V8tXjsF7m+uRmHyEBcbfPxX9oC5WzXFhnHb4Uipr+2lYReCEoM+
9QiDNZIaf1uZ+UHFkS0qh2ouBJHRRUbyAKrbUlAdQkF+AW3xK2/m6VUti9lN
5S+XipSyjWqLc+wuE+DCTkK8U6/bEo6WK613GShGpb+2kGyY345dc8S9WgJ+
h56rmL3u3EENyI6USpUMka0gOiSzypr++8PMKkD3ucev7+4wcJk0kJ4p96D3
4cuRq+inpimwgxhUoJZMEBvf9/m0tiNg37gZCQtOLrss6OUn0p7QJzulIA6t
Q/+IcxJEr6VGJEN0yTWmaN0XJ8aCsUX1/Mm/fKOD8EwUu0/1eRaqJ0GGidqi
oP1hOtDP5m4Efvr0k9PQsrZUVIKGAyZWkIn82eqRSk9b+ny1iFWhQQ55xHKX
/6nkGkQvXCogbOz1vgW6rabpDX/qXePFQ0XWauJnDEA1YIZgCeArpBZEFz7K
sFMOvai0gEpKKX7tDsnVmukQH6c1PdeX4Crxgj7zHcawesosnHOwn1yp9rmw
d68PHQ1hgDqEMKeGFuULPyBZgPQV0ucDym46CKFCA/cVTCquRosDfiUJOeVf
JTJh3gnRRVYrhxtGjAivGbkPp9+tvVZViai5Xg5NDaaZCdLKd5SSOcRpZctp
+m6mi+uKoNds0psUIwXERx3ng1VOXjtmBZYbgeis+5CeWI8wWCKh4MZRinPA
wahGa2BZYZhl9slzIhjsBFHTRwv7zn/BKxPnnzp0m87BeWjqRHqIOJ8OaafO
pmnoya2h/4URsw64YhU2+QvLxfVDz5ZyXLtOn/x+VThQ+LypHRrPdpZZMC0r
RxiRlyaSGjzlQHXsCFstKOpjimLuEsCLM70CIayJI1TwVpAElt32+weDG2AE
pdFsGMKBKQn2GboiD0jzMPplvRtPl4JBODa+04ABCMrr7EMYxfKPldnK0gsE
SWTI5b1tk+pDDfNYh07LNqysocTqkzVRFG9b/URi/mxDgasg12dbd02JVruI
8b3mc7xvVHq78f96Lkv3tBrGxR+xNqfbPBMiJZfi/NYBm7muA/KNEGrr1lmz
cGJHf0Bi4l2wBmV94gUFVqAvWZaZc9dQjGQLOaZqJqfUsNgiuBCK9H7m8On1
GansCtuwK8UyPvl9h7wX1L4jkiIpWOGrZAHMuPcaIu8JML5IDTRqQEtkRnRr
o9pfXkQFpS/NoRup6THDBmRVW9Tngx9PMX2+7ke15sj1nAdMtgkVhKUf3/Sf
x1A9kBckfAv1obV1CbvX/BUsKK3kCEeJbrbgnPxT2hrnSm/Yn6VgXvJPo6ZA
VFntDg0E57wKossRxoODl2fxekC5v6zMcNXxnEePSnmEgFXFDHbMqLlVN19L
ByNfNcyvFhqyzAoELHIgefPaHqsz4pSDySK4hFoF42Q+bMZpQzm1Sa411uq8
GDlFU5SSzh+W2hitvuso90f8NmEY1YLaU0YRJk/CGnrVJHWlnEsIvLok850g
7DjMRKHhzSfYtjuDXfMWsVpnTw9QZXESwvedYpfiWCjdBmStsw2O/JW4oPd1
kPDu3PK5yo7w3GfxhjALVH7urFDWzSPCc5q64Scbi/pM/md4KKo2P1cKhMQp
1J0srm7hVTBA8F/9YMxrVccH3HxiVKiR2rZHzvhOkYDXEgd2RqwIfwnsHcof
uMZvCe6FxpzhhQEV7fUxKm+yuWbgMMi2f7A1t479OsmQw+iWfinr6DeVpI2V
5lO+UZg7r3D+nNhiTeHlCdbmCA4SfwtO5D8INRZoERehtulf9srUwWUUlLw4
iRs6VAz/5OSZ23CkRjHA+1LwY0HfMfcngj4Mq75319d4d3TpWi0TWX4vr2e8
TN1aQKIl5oI94Wx2h06uRg2uEW3IKJz64tSyGjtGVp2tbAhtuWhPLYMkSkGg
NoZLeB3fXrXu+Nu2BUI/KnEyJy9zSZ8VjXjzYv9e6+caHGIonaZX0UutxfUH
ShpYHTCrsB2UGVva12vbUuuXVYNiI3oPP29az+qrC0Cp/bjX8CtOB6EXKJ7k
25I18ANsM6v5ow2UPSD6U7FwNB8wwYJdZdXZxv19f0jLkzO5ET672h4S2mmP
8Ta9iqiG5VhDuTxyCZQJbgByaCIFOgZkuQQclJforipRsAQBSF9Kh/RCb+vw
kJl1FK8gA1uztXP9fnWL1q/Us0IDeCnecUe2/WhVEccJn2wYSIZ7RIGMGDUX
ohikBKejiL9IYiHGnVXNP7BjNMbr2tT+FJPjKTSN+tLAEcf0nPzXT92e/2bB
kSaMYJ25HuRGfT+rdA7mI45W8D8VNpElLygt+9fEfUoM8VvIJ3xznyrkm//M
z583OS/8a/QLs8Rd1uFg1kiri6bjVSI06+pUp4Cwa/2GYmiSSgOx9Ndalc+O
in6f86BuJJCJdfB0aJtfRR+Ndre6VjrzGJPAwJu8wVq8/2LeOa6UlB0ZtZDg
tiJtmp+r5AEe3Xh3Op9PCgdTfM5wRWONHdf2scio/5BOg2z1dnvicgqUEEv2
b1jWX7TMAj3DbTOS+qhU4l+OwFK2b+GvXiGQA8oYjUJ3SwEpRfq5MFNpr94l
udA7DPj0Z00oPIPpWPYfnuyYYxgoOH6qk9SZ1mspzIT342UAnHjgZSrDi9ub
zkZ4BcIrMaM4lnWGOFEuh9kw0PFZGC0CFmbjR3ajRkEKfNrBtGPBN+cXqarG
rgmz4QxnNssJtlG59tgC6Ve3B7y3fKVg5SRkJXz/xIW8mehS3TSHP43Ji4Pc
Pa8snH715+u4yaKyDgIrK6jJdUA2qSeSD6eKIN+MRTyMymrZrQzCSnbEApLM
WaNamrlmxUmMstACAh5p0YJyLeSyMDqm7ZIyTBYlW3SK8Sh3+LdOlFIMAS/M
/fmRAQ+HgHHxu8cPI4XUeCOyV8xdSELuL2AQlKVUt5GCNM0bAPAkX3KQvUad
XwUq5jrOJ8Lz5MjNAwIF91ofUWI1YLcPbsK97V9D2ID1DB50UsaKJOLSz08H
58C0h0HMn7ZfwlxvuSgvahgCNRGi3EsxxJU7wHuiJgaIqcPkrnxZ8qdmN4NK
MtFoMMYWDmfbFV85bKU+ObLBAqMQP0NqYx3v4Py8jDLT0j8bYliHr17exMnO
rqxtBHDLuDh7rVe/ZIjPPqRstNFRsZq3GPsn3u6KyAqvGVPV1P1IHqR8RMO1
pBjNsoJXy8w1GXVnLZxbdfRySizCD9VuXyG3lrF3FpNI3lZDU7llDRVlDJMT
qmY7DqQiimC5toUn2khUnmBOnBAPRihKWSWS/kpdK0ANh85IhCl0aK6/abGN
EANOM4gbJf52woKHkLfmOjQ47dzg+2LsBNPXVQPGInlk49t9Xz/FVRR4bPD/
XKJnx12G3V3fRTpduiTna+8Nft7oFpBHAmZWdf9bxUe/nlRDgXajy9Vo0E5B
thoNuCygbN54494/UNFZqfEBw+lyVGFEMyla3gJL9F0dTYCYrZCbLDytO8k7
Ylpy5+OPt8bTCu+MMIj5pmPp0n04TYJ+a8uUjgU4VHuAUFnFmZJgbpWQzUDe
DRyZGarnQRMhzG0yRMwlyVIW7E4/PXoJPCI/nMXaKn+KuQXO5dutNGyJ8fwd
wTSpVM4Ks6M2Tv92jw8g3fl5xSjKBbPubQ+HJKyHVnKG0pvC0mO+gnmxSq+d
epO7VW712Au8Cm5rh6vNxH8dY3JCZ9SPMEwIVB9cwRd2NDvKaN8SH/++i3Pt
qCmTmPUvfl6rCN/Z3dJFHkdQeoRsi1qExTPYtPt8MNVOKmT0YOFWa0V5vS+d
oQ2/f8mAZ6cVMirNMfsx15UjypKIaWHt5VsUVU/B/Yi4KA08z+6M8vxmomsm
MHIVGyLDe8QnUr/WNEKJ/xEGd0ErPHYJVwjmJ+bQj+cqMc1/ujZp0AG55O+4
K51nblhowe1XV/ByjpBFTqpZJBK6AOgay4pF4AyhyLVjBh4j5sok59dLwErt
EdgF+sebynR6e7lo/sL8tShE4nxHr9ghxkbBcxBnxAyrJ0Xe8AmkvXLeV0BV
CEWodAOahoQ9Dfx4xxsSrjLxbN3JsWmgS0DrS9a41rPnP9imO0NHcT0fe11R
tL+fNsPqgy2P16ADdq5Yuiw0RpmMJ7/b3YEnDlyU6KcZQAWPeHv23lNVsziS
OebrRVeDE/y7cABAuaTNGmUQBoX1cQK5KrepIpZsMSWwXNUNqA86wrYoLGJt
jLFU+vPhSChtQ83L+PO2JJubMJcKTo9jalNbzOX/R3d5vHFJuSrPJtYem810
Tp2zHLt0tX8I4g4AKbopgcvY0BCKfY9+PWlrEOFqLlPHARS6a2P49ClEjrbT
3Ui6vcKfsJ/q/TLUrEi+hQqmnaJnTw8s0XaPMQZCK8PXjFa/BeaHTvPsrhop
6yt/txJpxb3+Wj4m3aseUvxPNXZSAIijdUMjO/bv5qd2G8pvFF/LE5ertZYq
F5lYp0U/ArybcjOOLxrb3l0O3ZBfk9Vy98LA/fBsvsnChMMW8Lw5hJvFctXD
m25VYzXRN/Kvzz10Kh8yFJsJ7Yxb84MkfGvJLCohS8qfzzbrOQLhgHmC6A1P
cXI1MyXUb3NdOjsyPaEphkkwW924sSAP4r6C7hCAQ2TaFsktiN+CVs4d/dVT
rQbrbSsw6IN4vkYMH/owz5PJI9+OJex2q4RtCbEpNtJtMPDwoREDV3GK/dps
bbc3T5GTYqoJPV1oWsJgUOmbKA1YyfGc5/7IthieKx/a5octim2io2DaUhTb
rComrC/+zSLWqAmCVgqqEwQJ1wXA108tCQtDorR6WRe6ynZkNTRCFmUW/ie6
3PaNQesttAfeujVyMN6x6wh/Abd/GjgF803pMh6ntxrseqCEMP/g0RfLMZm8
OZ8J5QQphnBXGsIY49/e6o8AXUIyBJjFHK0DW1F7xhL79ERs/73c6JDZF8Es
xeSw3U77A+a4lZzML/zNU3gh1gKpSb94AY1VFESuNAxWLsG1yVHKVnlq3E7e
uANfifTXAn0fGxPLAwZ0bh4a1ODdMiu465PcUknTL/jlI8RuMCP3IwfBm52b
EWASTBJddwQrZG8pRsNIy0MeGTtQ22tVr2R4UWKMYnBEFFNUgM4fFhnU5v6N
WBvqHIcRnOeCzVJn/YWGFBNiL6ZLDacLAyEokBy/Rwv55Qye7QM06g7KSuy6
YzicXTt/JXfFSNank2T9pH9M4kTjAYU0Q9Obisbi2fP9CF9SEmDsDzY1uNUa
+NU+wWGsYIDlvc+tFYC1lUE0NArp9RHd2LN+ZYTJuAOJp1gVbpvbM1jWHhkw
e/f7tsdnamDJh2lyr/ej5SqE7uCE8S3ozPEeFo/gthvFQtglTOgN/HT24J15
ccMBYhxX++9zEjoFenr2vjOU9+PIsr1jBn0yKXdpnhrHScIoSjimB2Ugkppd
sM/z2jfR/Bw8V9hhtg1o8UbfVJXrM31rpApviOh6V2pElFM6OzjaOFcLlBU6
KQGFx4bu6Kfcxz1H27R2qN9StAmz0cfqg4fhOYtF6W2wl3sHvpG5rPzI7YDv
XbNZMxcLeNDSAYIXa/6RykJA5MvPZXloxIFIv8ceAKlTjBM/GdM9QZUFXTKk
QjEheH7xo5GK/0pmH84f2lnFFn76rin250Tcxc/IPIAM12/dt7yzLlUvzolq
/e5jpJdxitLFD8JvPJGZ1Hdm8/wmUzqMeLXEyqjuleBI9Iprduaem3xhl54a
dRICRSv10+615jXA11TmyTElZqStlbRHCF+mDukwSn42sTYtPDx7JFzi4HC3
uAkjFTmEtazRtrAyfclvqr07rRMhaeMyaTotcTrxBzrP1MST2kNn/+/qvI3v
QVGKTynQffCrUUoiCZ+E9IvXNjXwlkVkVy1ATb7HbSHxTSLwaxiahXl2Bt0l
ltUlLZZ79nKWbriZkjppLmJmQrmNAoK1TIcYVv38SpXJqmyLNfDSOh2qKgVv
iemP8ph654X9armnwTre3h2w+ilhTMLk4ub857RF7X6ydRYCSNkP3CoH03Gx
yW09LzXICZCMmOFtskJzXSRs+SLVDB+NmO0IzNclFjvBCCuX1SAWAds2hUxE
UFFzS2hWSvHcVOBlDESHReJB2u9y4dF240Nor3Tz9dLEFXTb4nwF/I32OAca
OeCU660jUyTASIt9JhPd+SQtlTO6MwUMIBN3jhdV0haAe/CS99uvN/T9LpJk
kT0yF4BcjyxP61zNd3KE5U0oAdwxSVhaqSuhDCSczjeRjh0ogTjWyzn4pbIU
gXsXTUcwlHNRdCbYyvGVbyXO/8zvpoDkKQnWn27T+SrqbiaryHv9I2HpEUv9
f8B31JpVXAn2Jepdekh9VJj1H39J166WXnRwFvgvewR/+1Ar5rGrr8vKBcoJ
vk6n4FlQBwM+mwPRXGq5zbCpQelOnN2qXkRZzqLF26cs8X/dElpiSfWV0wRT
h6jVorkSp7vWlezRDXur3Fb3yfs6TEGsxBoe9Ks41mUoIoJ4+wSvqPVtKexQ
sZdo7mODvPWKawzqwbTyFS97384sphRZ5gxNFfC28tu/eN/NlkeVGrOid06l
ZiemEtyqENLc/NY8h73TsGDYgh43nh3HSM8UTaZgrro+OELRFya6xZCRQERU
ZwzXALtOlkeFBmpzeFxgMaqusTNhJsrtGZjwtx0vRSxenWNPQ68Oaeyuk0m6
aHgaqaya5ff82wkinfImc0QJWYArGIyTJoWXMzrmQr/uMKDbhuxzdP6xdR0k
yLaz6/ENC3TlhVYQp8txV/L8oZBLK2fCWpi3fGL+Sj8qI8UEEP28Ods46oym
bkdkm/ulDGqCdMGCFxaWKyVult5wCQNoJWlDqnha1N5DiXRpCAhgwWOM52Uc
GTvvw9O/xG/57K9n87GqpGvmDYfw6nyxvjM3kZ3rVSX22aGoEvzmXQNkTjlq
rZBobi3Qc92gXZSjZiI7T+tEQgvpzdskPV9I51BNSZPQgMiBOpRyqkhTFhD4
1mI9pPcykqzEBcg9fzM8F+NZyxAzUOqYGQm1X0+vyrCPcJtJUsncwxau+8s5
WpUhfK0zUutvX+VHErJ0xbqPn22aaqpRkJAdhFArOkn33b2aVu15c7NXowo1
VrGYl2ysICmg1dOyD0x+jIbpaRedTzto7wFhDo0v0mCt18cye/JQTm8woRtg
kJv4NgIKbT5mTfJXzluz0s/F3eAdC3/tszk8gWpU8m8sgD2gvAxvYicBrtkE
kyBLW8HT7WkVcd+938ENXTxfRxkHoNQmK8r7/XxodGrM3Uivi9Phn8+ae1OZ
8D7MqLkQ0O/3Q7AO7ztExo071akyLFOCDtEgrSRZmPS/3oPnUzmBZtsl3PgA
m0IHj5tf3dtWMYpYaHEV8bAis9lZrloOwsFtWVCwoWVcepKwQZKZxkkB4nGN
+ZJQqQifG8g9rCMf1ity+4lLfECqov7BoH1nOpdFLKEOvp1pnpx9z7knGffp
VQv4AWziX+MTDBMQvn7M0/2mOx7PFxq/1izaPSftZkNlBNYdYbbJ4OTAdyo1
EC24i6e3iVUx38OZrxzW+pAvLlO9Mi88FReAs48x8+9tRQBHKsC5aanioq5L
7WziFGxyZc3632barldommJg+4msTGTIh8dLuWfbvfKp2dnqcsiAzVUS8J6u
G8D8nAYwJxll8bYHMQjgZX7WUmpQdwN9z05rKdgJYqIpqNqKVE9okGeebY1v
YgkgPap0pAcfm32PpcvKHZkwiojuaH2hJQiOT0KL1Mjb+X6p74jjhlQPRA5V
qui3RMc92YKq9baq5xdZyeaeeUstJ4XYIwi3zUBNCUfDF3Vg+LRzPCGdrbkl
OHrJn817/if5dMPL3KGKCycLi3cFDLy8+zuNLFHj8t7s2QTVOpOQx+BMZZtv
ozI1QOGTpw+y8g7RX6cs241rxQnng5PM0rO8KPbPGjhhoG+ovzgHP9pg4VX8
9BAoY0gcuIdbbMzSO93cmDrBorfRNEYJZrCxxna3dilo76UXnnmu8vglf4Zl
dYg3ohygrrBy+lBwuFb5kv+PYDGp0FNIk8vroETQ3bfQ3fYB31i5zj576Wxm
1KdG2iLfvoZBYll1FHBXjdDyuyoEpjE0ZS3GGsSX2dNKNn/xTfBSltFrG1/z
v7MjgUH1uLuTXUZNR5H34dl25TjxKSCW6zD0Frr0o5qaGT3tO37wErGx2mfn
lyJ4RCe2nF0f6kPBTWt45XWmGptxNxk5bHK1/Ni5eWiz5J8NWNFalQE7icC1
uVA9ousl0z9l/3F89O4IRxIMgYYWdDphqkr8b/ZyB80i3vwgUwAFgl+fjlgL
nc7XSex4JUAqGmQzkTitQY+OkMqxz2Lcb2qCLA8Fs2d8+VV8uQS3PxZ5Rnik
HNQUprhtoPLPiJ8VuiApWTEtY+HazD28vgAlphUCnbCGZk608KpKi7WodkV0
Vb+SDUduowm1pfoo+4miQTaqZHmCyRhGbJXh2cvbgJfJQSPSwUKvXJGW1ZMs
0h0Knzwy6f5UXSfx7dtk41IIQUS0v5UHJxEf4GwMQj4lAZkflh43SW41coSp
9V8AC0Qr898CnzU3xYsnuPZsNvLC5c57JKL0af+6TaSfqvd5JRmWi757zfyY
w1VaO9T8E5ytyDjaTvmxZwnYg8EpSdswtLMsE/+tut6NfXagxgXLYCj7hTW7
GblU3yBzzqLZUHD8bzrO2lAw2pnwQ5ZSYKS7szxdNF4XqBeRftPfhDdjHThQ
MYWJAWibHv+bWs674gemFa5UxkhzNc3HPV2tD6x77OTIRm+JnVkyCbGFkgS/
NxEefH3id/NnquY7VBA1QOF/tCuXDViXGXjHZQiAMUfnNIup4xauh8CmhTK6
OwBcpQlZqrZ7tTLBMGg6gzJwIkR0qXo80u+7n4HoLUUx+Nlg7JJcq//dzVf8
0QRBMXM1QEAlGdH6XDea4Am52J22hXAf9rLtkbUaCl0ShGhWDNw/QIG00d2L
GOZEoj4gyvSogDw+pdUXs4+8XEaxHIf0a/yUtdLvnG/2RK/ILOZ1n9JZczj/
b1o/yKp/TFcU4PUzDbDXfZ/PpQA/Nc4DxmdAh7iw2x+YmAzj3Dlio6h+A1FH
GzHZoo0XMydPhSQVbVAkPTYEluWwO7nd/Uc2uMoJp50JwaOwXhViACht5jFd
4tLoCEi2jdCgLIYqfPWCFkP8u2QncAroXmyLU34najgyI7GJ7amjpb9f0OZw
pjH1g9qwxNLbA/jdUO5E6HL/wsohb0od0h8hVOS+Ur9whAJoxK8U+igzioFT
dwNlS9FSkIt0dJcauyyKuTx4rH3SEnUgvzDmYzd59VqsKYxCU0myPgMb2o7P
kFjqD14xS3dr3sfOdVYF5LDlPOPr1cwV0oppg4J+1qRLW14XjXiLyjmCAHIM
wifEJ+tSfsHo2mLTCNLFjNb9tB1y4KcOn5fqwqbc85bYNl5oTEfI0bYUqOAX
Dd93mFMGwnv0+vrDBE53nUGT9bHduILxcBsJmx2jhjZLyFKFj0m3YLjOp/nY
RvPerq41oMk4w8dxUEe68W+dztg4Ky3vNbD1laWT5+vn9en9w9fzzt4D/KUb
gpZnTJvw240zIF/oNRfTXiR4ljyeZltMrjzGSUHxVQBdBEWaAnrPgb/WitUT
cVhv0iyn7nILEmA2jFCpmuuY6cTp22N8RH3+f26olEQRBgROmDa8QTV+X4m3
9aJGzYQcFFOV6GJoYpg7SsskArSFWeFpjd8Kqvhk+0BLrQN+9UllzsXQN5zR
nO185E1k8q6mz809IiwVyi7Jio9vg2eGQ0DwMAO1ZyT18ppmbvAfrsbBYkjQ
DdMEPak8OeDSTU7Z5Pjelsb6Ipei6MpMBF4PpYvGZI5/lIaynRK8PyDQYthW
pB1YEFd/9zMv7nv0PrWrR/ogv97nCF5ab0yCxcWH35X2Jd68E/YbDsX0+Ij4
fGBxzPjAIWOgkbCl3Jyt0meWrF9zhMIBZeEBkASHDlEfiqB2dOV/cxnwKs/r
DO5GuY0YatyVmE6tYcw4JIUgSTSfmJjW1WTXSDGyIjUDZVgUCTWcEGSs1UIT
R5zDtS31UmHH//StkcDQT8d0+yuUsaHZZplwA2PZFSUgxsupeGaUkdSVavv7
FvkqY+1jRcgfjozZ73K53Xx+AJMXoFRDNi0tyRmR6kTXy8s6zHMjnRE86vwA
4qMmt6U8LgDK99+fvraBsWP1YhypRI35XGVCajJoGcaaqo/0BsMxMfBUu5Df
d1qUfgjHm5B0zug9DGjgVvSWt8xdFN9F6bC1nY/KuDOHRI+PW8s75XL3gFhx
W0korJJgP9hAaUaNjOTp+0P2ecahlwcSzEj/EmrqtEZOAAqHkKswmFBeeTy6
0erFnAqjT3HP7MFBgcArOJxpi6EK6IEI+lU3dCnMz1ZWfJ6ToMYP6J7o2Fu9
YjwvcDsb9VJp4ua4PgGk/NTiiceDNoRw/ZPTIh23L+GW/5boBBtIlszXcg2J
Mclahb0HQ8kQMrSHeigEfeyV5P9ycdo5oKZ28p57JZPIYDIWn2/B8QHPcnCj
p4KfbB9Y9RZSDEo5+3oSZzL26RjjtKyzA2zoB9szEzYRQ1+KfMTepObmbiBz
khAOGvKE+s1eRAjkXRjfY7Nc1QnuFchEWEFzQIrGAHLlJzBMhKgIH9qJsG/p
0l7fMMiqZZH7rzVytVgxZeT/+1GL2jUuOc4eOVYH6RG6U7emPIjxHA56fBGa
qWeLjHuAB92yZO/HE3OGOrl3e7wnTCXfCPOiCPV1TSvZQ8Bc4i7cz4U4nhsR
IRJnpez2AQDcjwn9GCDHnVDR3pUs9BEKE1oxnW/SS0JAcJxLAR62T71fe6Zz
X2ShgW9TRkhkCepp/tMfsM/AJRP5lihbKamsgxXc50QeSuCetJXLXBQ0KdOT
PoJUICdoSX6gL6JwPTB5K3UpuG4Wq7qUQNO9FQ2IXJ7a8FXVW8SESd933mGM
HPHOU7pP5ViUoBwVhl7qzVpSJpBHUwivkWOthcT2BXPavtP0CHyFcPKlkcPF
pYyN/Ej5uJCFoUPV+Ez4aJ3W1rh6uOJ7w6HWaQHbIM+E0qoBvOTLvCZVobTS
3ok52NnRHax9h0dy78knYMXec1K3ZjDCiJ9s3QcMUhCXY7C26nPnELCn3p4P
5AZVnn8fzf+ltG0V8I7Q7uKyKVBaK1+gZ5HxZXZ2scu9YILJ5qceP+kqi/0K
kS587NMYoHYXvOUg1EK05sYsJIArnVMkPSrQxi8zjqETaEMHn9yXQLNQ28Au
qhUJHCLEup3I7/zqrs2pc/Q97QNeWeIi0P5lzCR5+kM/mWiIFRpZCmBpiMrs
5umDJbF9tFEOv72+ltCnCE3n+LEyEwP1PdmuBC2S1WGm7mDVXofzqw6uiIf2
hrYqtMKn+c6PZTrryqIaWa/JE6L5h4XFPSVi1z0+S5TKVExqnejAROqIsMR+
Cqcr1rd6tGRDwNs7jx6nISkc3ykBSf7XmnzKKK0gYZqbeCqsitEPRDQXYLhz
8/q+DThDejxSZKU75mhwjvrEjGB+DweSTTwNwEUU3ho20EDB0Cma6jlwP5qk
ptQb88lNC9Xy6A4aw9Dfhj5iTdFaOclDsUotjSKVZrK5HNHsK9difKzC1oWO
3FCRwv9Wqlx3tyNVo8sij7xJD2SbwQs0n8OOWBvJwu1Hor4nLsa9XsqivctZ
u13aUnvvCazWXQ7gNoYanVLnJaWVE5x5ELtH7Q55MfKYc4C6EzoK2dXjYApw
TPVYaFSa1BwWlC+Jc/I/jBY6Dae8611VSu0UiAS/nwYUootWa9Zzm7iVmzXC
vddVYTTcfl3d7B9W+4fcN9e8aH0NdhAeu+QCRQjk9ITBZ8RT9ck3u595JQrr
9YXC6I7sOaFnMuRKvNG/ik00SGOWGuCzic538oX5fTjn6mqXv2aTEAjs4qIH
gp4ESESla8DYs7qKh9eOc7+DfFnwHzDYJyhr8rmEDLMbhfLldns0BOw4PUlt
W3TM4AIuxIgBUdlf6JYl+oFBEf8kWZM9/q7A3VEXNlAhRqSm2s86H7bN2O4H
1rpyt/UHihgYP34gHtZrb6dOEDeMDjuH2/ZmdH1HXh/hdItgiZelRMOb94W8
c8U+myiqs1Z5gjfmI0q/t++2Sw7KZZ0DzyzsodV2wzEveTvnDvuGlKQkh79w
5AHyPocepzx1/leJbYFs9vtKhtOQk5Ey5Nwfl2X/IEybCmCxzyC5e55ADWxZ
TW6Rl/kTgb6crJodMJgYFbg2LCtImQ33daOFPSUbpwyzAcmbCDW9JNtBS21a
I9EnIcnDY3l9TFea/QwDQZJRWCiZKA2WSSCGpiiVcBiderDtYPKfsppZAzhN
Jhh9wmCnYGissbYSZstuHXdnfDheviz03VWmwCDtZQrGhqXUSS0VdEMVUrSB
gCDjlRRX/+pAfMp//obpyidjYmsYJilZRohoqYmh9HeOnRYAo/O/1RYhYiWx
KadrTzb2PcYfg0Au0CMn5PCjw+dE0WW1aEL55l/4XBiNveH41YXaxJBmkT8T
dVRgiuNGcQVxwM44LGqw7ADULpbyAB86RWJtEJJy3kKcPsSYDTX44JlG4Q33
rdGE4LQabGfAjm2P8whPAyfaQXqz2MOBklnwYQPThzqCYK2PE79cUGywwC5a
lKkAdiLP71noQJD5d9RC4wBN9kVYYtcWl2vhqL+vzn0L1UNlOsA/6O0XbceI
RZqziJvHbe3EiPNZm5gpKty/LWa4eVqiVYrSu2UUFMRzQKv51KdauGdN2TQX
gC6up/haqb9bkh5wohqBsJj3uJton0SLi3w65Zl1kx94FhYvEfoBaEDj42Oe
4hzo04SExKs+azPfKwwYuYR2okP6AYH2aBcDG/3y4gIXDJlrFlFl54RBnK9R
5uAad3O1buBqOhadKCwTzy3dJYUEUcbKW8m14UetndzhPgtQuVCWQGdkdzel
8bf1l2fHaSehhqoZdOAaf++dEEbO7LRIVL54P3qymnQCjsgtvhQ3o6UsePJ4
kGCiyWCJNH1SihbO8AhxV/4Yc258LlXf37/J2db8Lzv8YphiNy/DkjdwDzeZ
HQf0/AvFODsELw9EEXc9CSvv+qCXRRCtQr2Xgxg55DXGkuXGhZHlPdRRljdY
J5nbPOFwd2INK5AfnPUpCNmTM5VCfrFsm/qr2DtiJyFBO+9zjFDE4n20ImIY
0VQAbuHenP750FRIEucnVTDS8/Vh2FoKWKJzYnU/kys34WKsdATHfkVrHUbz
zpa4rYkPU/vikkzbS3r6GfGBIuO+ZTjM8AAIA04Z9OgfnKH8rVo0UiS281+R
dtL+d5zeIwqfikwgnqlHEF74y4jToOEZgwTDoL8PrXsQYfGidBV5pRwsO/pN
F/m3i84d8JL3WN4OORbQKFEsPRujhK8Vc2QiUcf+PMUAHaPymdbdr15MpaAh
9PYN5vkk5IjObLADOxsnYdcEYrx41rnZmhcivI8feSsAfog0AIZTfDYiLZKW
iYL8UZ1EUWj0IvBBb7hfbOSzl7fG5tLtDz5TFwm274JdPPnSwqS1Er8h8LJP
1OzhXF89iEsnKnXCFI9VwKYZ/7TCCKK2hi8/0ZO9FtcpimjQyXiTe/xcpvj+
MVan02woE5c6Orh+UJxrmU5Ndlz6x6Lnn8T4LH1jIkrcgUS/1VHAGAzP3DXz
3RRcZlYWGmzK76brN9UoHZDhtyS12LLXgfvMP5I7DSFONURfL+vXPsNRyU1d
kK4cvcb2IlOSZ5hVJUW5vL0PRf1MN0mDUSgTXeI3NHqNwYJysHU2qnpuklG2
s9Aqe0jtv1+utob00GH8Ir76/bzVM0I5rui3yEoOxAav6UzS0iDS/sRa6d3U
kOIu5ZrwFwCILwnO10kdphqeWuAsCbVx0kUFnr7Zi2q4hpO/Zh5/pqUsjgjp
UR9W4tGFL4N24WV5Ss3PXwh4IHQmaQV3vjH/Km+8NOoXJ8Kwg/TApE4Kwa90
16iUrqF4qkecBo3FjTcIkOWEEUbvTZqLhT8ur7MvHF7XkawpgcoNVgv2yyX+
PfKQa6wO0VJFhd/aHur1LKmWmlIrhHh+SxTIgjhBGJ5VzgH4BGMChOWwna42
ZcOdosUAZCa7lzqDIBBJTnphddazDY7rRmd1fkSdbp1XQQO9u059+Dz8QVdk
ywWghnI6ykHrgMNiIBFfIY8VLr63sHw2DogwJWxglTTR+pB5QwdLL1vXXqaY
qEwkkEXFVj3yWGmXagnRnCDrs+vQ2143Gctl2tQ0oAA2Y3fmy/mBPguc3RMa
klUI89lzJQu3qaCt4DREe/wiXrcSUWIbG6n9NfnpvWrLfX0BKxc71JjIjrsf
HtRQt2TbOGKl8O9HzK55oPYSlHWFoIG93It0Fzry+c/Sf7HX3/37g702cgFX
vjVQ+53QiHcnNYz32T9kVui3QzhIwqIYGxiZxXNBys0kw5/tDbLBiKYhUMUk
FAzd3WVD06V4bDt+Tuqa0oz+sOUn4X3CVccQSL6dn4yHxeDLV8eRm00peZUE
0/Vzd2178HWM0dPXB01EuIxXBTcHJdw7s5y4K+JZR5bM9+5CqJb6aGxMvSLi
oJHnPB5j4oj51BA5MDzXRQKysCx7pmNGEDalgi0a5l/ZDMecpydR8BLMWs3J
cBvQqvH/rY+M8itKD5iaF1+0f++tm3puLV9yxZVP+6Wi+BgkNGlrmfQ2uBqq
DGRL0iu9NX1mR2k9CR7jVK8V0kgeQxRGkam/jVqlddTDizo6TFvtMFoGmdPS
bH5cDCHT+QuITpwYxHxeOlAK0MihgksGSE4i+BJWExpz4H9y3I9yAd3Re6ue
inh1bce0WDRS2yU5xBZ1iWm5zTtHDXfEIX0D4rT5ZdAerQqRI34JlW9RwWGd
S8fHLghadjpNvb5jXYIccnFaLZml7L89FkLEZ0+/U9ipQ6qZTVQ1LdSOeaMO
eQycCn1m0UZxoHNa1s+BliBdl7B8cKQrIi8wIGBeHuTl9k0JcJCpqrXYzVOS
0v7aLr2S+2kYW7AnU3SkqYDA4/md629yoRiRh1QCM/x3K3HOjNqVI4g3VzmE
Om2b7HkBDeCG69cRy8IdmdeIGFhp4Vf3h4YfSEoeyTQtyYBQTKCqTLv9WcPC
Fyv6e3tQ9MBavfPI0ff7fmEr2nsp6OjKRW4YnxX7ry4GViBGq1j10RFrXq4t
t4fQhxEPzDIbium13rxoZ3GgEWoFXboVB9boFjJEJt2h+17C51Q1HQMQrecO
tGCu6QU0tbvDnBovPENQageQfEB2CvRqOJ9p7AGytwYOUtCnr3ZxMYjdbmO8
i9agrmomXbPZqFkEFZIE9WcVT/GMRfmBhnaxHFWWmQac6v9zZLxKZU/TWOCm
JcJFMzi2PHAHmFG5jfWlq4RmvF4bYEJiZAE+ujOJIuHdjRmH0ZLSGZL+TTRS
kJymhn3JDuqibKXV2EXnD+FXvCAHjgk4yjFYRWMZZiBrsKwW+PGXVNDb6OkE
xxoP/TVvekGcB8SIgNTD6lPhUDudqNWayEdDCRH+FBihUQx4Ib8kCfbJSp2r
SMOlBro9AjHKAOwID0oVA2qRLfoyk1/u0VgtzVupo4QnV3tM3x2Qc4KJQeDk
goMVa2J/5c7pY+g0BlfBH6hBGYi7M2cNMaL/akw38WcxjhOaC/ABe9eu4si+
c8dq5zfsDjdBv50D0jwy1ajmm9xFlvjw5Px6StGr+wP+ACC7Nm7kiDBIOE7J
nOSVn/NzjyD3nSYJpue4+LabReieiNQI33iltQp58v0LTzIkbLuW8/T4420+
Kr9wgdP0rkNPeYkwazXk8GPAKHGF2fP5CeE2Hf172REK40f6gJNs/h/ip1Md
cR4kQpblernCI1Up9jyYJWFPngS9HP10pX6Nln1PxYF8JFyr8wzFG36XV42S
bL5eXAZlrVTV6O0RBO6/3Sr6m7O3gLQVgPtBw1il1ZUoEeAPQjFL8j/hk72m
vLqNfnwSfBkWjtZcyEQp0r8/1OErUksXXBAzstJcH+DfJlslRbLp2fAHP2o2
as8bi8mwsh1csooeIOkcUQFpuKT+FjmH7qg0fqnL/40Th2rtzozXQ5o+SvE4
KDT5YiKlCt49QWh+oSVvjezLv0ik++YKmWGr6egxqgeVK9T96tUi2FWfbxCI
PQVR6/UdJ/g2aXUfyQnDyarNMDcVNKC/vPG+r+y4NxzKRFyiEBFK/TwIKKpS
P1OvJzLcFbMQGSc41ziEKhluEw2jRSVhNi0Xb8rGWa1MLSGHxfSlO1dbzwwp
QzBzKqpC/0SqQIs1r5wK3jIOcUafPBF7w8vXxWFt/XFCEy/Gi+QFh2n2AMU2
no+oaf8B2Q6TFQvww1Hsayj/GziYjd9byioUFpDuHsjWd6sXyoyKzzJSGdwI
1G2Q2qjhCNPmowcnt4WP55gFK5q4W/ksbGJcb2DM3lk0IBCVyL3zVkiVecjN
dLPiTIMhWcC3PKUYUpdDWVhywheznED84n3HKwXUjWCXyZUzwy/0AC4XZoot
8xZuYQFp2Jg086xN8YcUivrwxQv+n3TcZ97/d3KhAoIyDt2WRgoXUb/u3lZk
sNoFyJorQtmQirqtcE3YPpjggXfCht9YfL3vRATJSRipzljt7zkM/i3MreMb
J6jhcV754TL9zZ1wocZ1JLJei58SPp7X

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe76wdOtqPzYxbhxEpueQaR7D1eergdxrDN6X9iqtUTsM42FgxnD2kGUIELMVzFVyGViRSJmFGJNl1broZ7CGIoZtSKoqV19c2s9Sn5zRIAI7fgXOp/nekBWPyJ4H2qvQqKQPAKctuCs1VEZ1lvdcGSauRG5Gvl/jibjJ7OXpWKIxdLkHkMLWaoGvsF+WYaFIa887ihgEF8rpbn7b9F3jpx/9QSKdodIWUi2FS3y0z1jPekCxIZ7dAPvXlcRevBA/B01aeK1OZe6fpMYWO0QhavYJe+wFEDxb+ZHCFWfK3Vu5lBhcRQkw+U0h870TmBVr/yhwmU1C9nLS3B/eR1lInj3lu428jFYWx9IT88x+AJ6g7TT7/wKwQsohULyoLxIHzfW4WyfqFfLmyLHPt8X3GeHOGqlK9y5Ps1zqIaTtpchk1Fo9jFfdbNrDcuLcLMfw/ABY6t4/emDwKIaVhtQZzJxonvlRKH+J8frGSHYnO6H9FSkrSK9P9A0A+mY0ZfhQMdemGMMNZt8suuwSZWVl7LSnYI9tiYx0tdJszACACu65oSGeBeD/BLNdmeVnDXtQPqtTU6N7Hg+xWwbnH7+Sc1Na6+L63YwLYgnox2SYzhiwCNCtsFpvSHLtqUOog1QY9/KrT/YiQFNDyMw/wXugCLFRxl4U2pvrZMiHYYEY/FDOrLEI4+Y9TAx2CWesQE6bOy3GuloswKHty6DCF+bF16YakSjXybJ0BM9X5hNgaDWWG4Fr3Us/PoFr3WFeDP4U6X6+bchwiUhHt/teWDfs+rKS"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qPpcjz0LslTT/369Mbwr6IQy4MsWm0o/p+BhHtod3IjCrEQVSrQ2O4Qfql61
tNWxlNVhI30f8A5qd8cAdXWajiGd9QIb7wLDF9t5a6t9DuDXQEV/AKcytcnq
hAKXolttzp5uCKHZ9t4wsl5AWUxKsKOrVasWkFszj8h9ZNB3aaHBqvvrnv5g
PYgLxBJG6kehp0W9YjrkGWZkNaBNZbff5LLfHoqQ6jL22o7B8DEMF7QRlR10
7XUIaOTRy0E2zaXFfyjXiQxuZLx5oM/4g2tyyqND62To8cR1MpG1Id+VARzg
zBWieley508qxY31+WWYqdoDY7DKo3KbU91KYp+krQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OZrvK7oZqWuMxF3z/QK40klvv1KFj7cmzhkdR6cfNP1BAsh8mUNcwQGHLbIt
yPCfr0TAE6r7/hctKqdiwc9TjJ1NRXT06RT/WezVEqsaCxHXsjQ6yc1OC7Hd
XPDmi3BdwVu2oLzuTVd8b0qu2D0NZgqu3F3od9tkX1c4zxAM0kuz0MUZja6L
eG0QP6Xp2xSssxXM03AT7DUnAn7W+oFs9tA/n/Ezfg6VCrVOAnxscnqg/hFo
RAiFmbQSdxVyhucmdIy6YZdPaKyLjWkFY7LYJIS+hOFnM9NEyIgu5p29j1Nb
0xr1n3IlfuxlSAYDVPwSTyabBFfHzMBfoPfbx7J25w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D/6mpqF35ZyWh19SD0f8A/X+n/l67N9Yh9LHxUzwXf2AwskN0BcBrURxM9Pt
FAM5KD/7OnQz6h9G/tx10nzTSLI+NU6gt7MB/Tu/kICKAYovmJl+jwBzJMl5
/cEbFccxIVBp3NokyqWj3BTp8od1Mdfvbl+VaCrLV0Fxi0UfE34T1ey6nDxG
ZYQ/HdGNUhkt9jZQWJdQSDgIZa6picbn78FwLGsRuXCzgfl63kFWnmTw/Abx
cViAaXeq8plrplqpHADICLOGaEWshFRJb6hU1XcYuufICEo/1ixcruIPqjA4
GyOR8Y7UKl9OBNyY2YQRtcxkhPGhb0sdeJkg1+sWNA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nXlo3mgT58rd0yqowiDIsyLNGEA3BBX8C1eXmLfDj/AMXawW9Ju5DQj5YnZK
C+9wePLKPzjE3yym0YRTookwnw3rRAbbBzksjObHohjSNmv/jwvZZ4Bhsq8L
YC43lXrybtqOMRi/BN1yuM3joqh/hL23WJqbuAhblBsDkKUR4MaluZtii+bV
eRRpnbTumsF6XQGGR83rZ4dBItrDj9V4BQ0r9HSNJ2ZyuxMI8a6BkWIb/k8I
zy82YOZZig4lp339WUh+/9w4A+Njs1kjqgOqTBi2CjOtneTtXWwxeGkJrkGQ
bUp6p19D38/nOkKSP6AMSh1fbwMv9KDakmBFUA1Tjg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oktPb7ZVQDYp8BJmTiwNnx6Gb0EEO/zzTaNRb4XzVyQg5kAVykwMVJV2fu+7
MigRe/ElkVt3j71mjGEUK7SPddbppTayYhtff+kcIRXHnb0R8P7oytMdskWW
G5R7wXWSR0d5qO5mEItM0UrgknH/ytESMJKmlg04t0MCDnRaYI8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IDrha4+dQWSmuSr/NVFpW5gkv/I9hfdo3kwrmCyMuzXLM86YCf5gOsy+en2Y
qvQUUg1Bh+XEaGl2bi7CE4LB4C/ppWimHcCMXLRb/T1g8ko2BGcXls00yClk
vcSr6vjE6kvKaQdEnQR4fxCaC4J9ufFSTmaVnT00OZlF/ZTWQW9j0PVAeT5D
QwTZ+qV6qdv6u0SLvDK8qXPM+dJyPHeQ/m61UoclqGwpJBu5ksfSUHO5viO+
nLWXOOS/W3UwfTED69IJfmd9WSn/Tq0231glaTTvB+KeVxeB+krQg4Bv5gsr
i0OV9inn1L0Vj6k4uX311ybCw3pNchMKgSD/HQz0k4DGyitR3lu/rLUU/TS1
28rwQkSpaSofELhyJPJBT7sgJt55jeyRS/B98zvyixf55Mh/672sR33v+wH4
C0zdpG5P+S7g0kxDLDc0fzA2nS2XTNX6VM3O3ouIZMUW05oEhjYWhlvpTP5M
FEKLvxP3W2JQMZ2kfCnzEiVvDm7rWsek


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fzb1R3IpJtlOJaZEsNBjmFjdIGI7U+4/UX2uz5o06aRKqulp3xdNU2NgDvmi
RZQcbkRew4zNFmY1GVpVk1kspbZvj5Tla324KR0p8a0hna0OJltnwr9O00VO
RMVU3ooLpWWAmzjHXPMSfoVEqLKXWkoAzFzorh7Pct/5d6OMtfQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ioh/aZMSHJXmnRY2YZyWLBgGqKgkXqMtniuyrC9Y7JkBiyGQaxZvrtCKqPIH
VBoREetkMFEuqOd1UtB2LbjtPIjY4JQS5Ohk1OGvcmXNvOOMGKm36KyKKTrv
t+K79AVkXdRfrxftp1e9obZxCB1xOFBU9kXk5Y1b/f2LhPcviXY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1232)
`pragma protect data_block
I00CTJpFvLrHkFRE2wGEIMrdpnIRmYS5+3QOr5i/oqx6Rc5JlUdPPepzehHt
0WopKMIHYAMr3wIVxMX3RHVH3IwbLgpMYyC3gIo2crcFWkvFaIUM08GCSvbd
Ai4Ydj1t4npw0aeWGeHVWIiv5FzM/hLpuYSL0OcRfP4AogJxNf24pIvJtMJH
gY08gao1XMDSXtCxhBsCbsMrv8PT6CfmMoYSEkj+OjevSO/h+cYUJw9eJcaf
8KiuutlCGyQxH5J5TXec/xNKUGkfePrw/8kd3EQXFjQVYrvQ92F8c4/+xE1f
FLNuJ2xmxAtQfukSFNu+EFsVIbffu0Xp3AqmGTxgUDzZzFzumug1WGS1QM/P
RlrHe9TA99KK9NFQLPaGmE0aXxoiYVQCtopMH/P51TfE74SXFGl+bI0egVxD
L3C7cXP2H82Rfvxu9SKMQ4jUzkcz2EqcknxOI9F6SxhYs4UiFel5UKylo968
P4jJJ0VoUA6u7fZoAhBqG6/On930bIHLh5rPlg5OzXlvxsz6HpW4KBTtGaJr
2+aHL8KPvPppQBosSZaahS3X+jVbxKn85L5bZu2HhFqMwF8b7SX2u0dMJkEI
FWyte/KNKkfqsS+FUb6pH8uEvJYfyA/E4tpY7uHnq2xCnGk1CeZecV2dHtJd
OUisETYj0Bmimo3e2HaCx32sA4c8/JhADnWjkEYZApN+1KX8KO2wN9xfCnZ0
t6B7dYeumHeVKkBjRbDkYMYXhZf/3UGT+bkteCAsZl8l1naIF7zsNbRhNpKl
YNQiL0qyciw3KjGvPrz/N85z/uUKvqijYkdMkK2INYF6L/QDw/pio4GJ6kQQ
CLUPahaQQtUyPqIdM8vURRIfw6StgOVj7o7GVJaiJ98mFSxhwUeDeEy5SZzw
2Kc9O1RTG8uRN8Bv9pY264FsIf6XZZGzTzHFU75bTBKMtOMRD2fPRUK9/LUe
yJdjLdbXnjNUUHk5JT/SvfkAXvUeU6tcbrHaMz1o93rX/J7lIL65Ea+5tJ0X
p1rTMBI9WxmR76SMIqQboTgP7zAbj67Aee0RkNea6iATv60vcDZ1CZAuObZl
gOHLW7lBBisgVWLe9np0QpT10EhTOByr3EsaKqAYnwS7mdEjizC8tJXgSRFW
6oCdP0fNOK2ul4h212Fm7Y0OHNNM9JgBzH1grNvbq29cerPCIWYOMaIx2lhF
JMHAzvi2DP61C4l66tLgy6VfoEfqOcqjYBsaj9B5Q01Qr1+QmSO2qrcnGnC6
Kpze6hCNvKXl0Pl98xY2z30WuRm/k1a7nVD4TcdoMH4Nqz7sDAn2Zkz0zENv
my6Em8Ttnz5+uckUd1Nc5JK8BAbbs6zq6x3z8KZuQ8MYjqRVi9o6oVSivN3T
kQsLu1VsVQ9BZ0CjgU6a1/ZlM5HCh6iEVC6DBJm/TiukbupkPoAvCQT+OMxg
yylPoQwTj0c5fm4aTkCqO8qYMPwblH1sJ/Ap86mXfdKq+HU0EH8f+qhZL6En
qD55JZZfC24j7PgAOuA8Nkneh1iB/RCLfmLlsZIfnyZVkf53F9Fi/WiRfsWk
1pLZnVIkClHCCvSn2SVzuX9CAgtkU/YIH1hbNEZq4+cmIOF8IOLin0EDqcmk
E+SuWN44bM58yV3F6DicK7g=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI28d8wF0ItTR/iDdk09cSQSqOeLM3Owmf79wQpnUemnVeHoNvJi1TKRJ9XcrvQyU99hk+pgKqbZ06xkS9JUIQdJSsgblCEqXhDuXbOtdYv98vVpEFCp5PQFgWLGRFz9mugoi3stBAwSltu0fccTqCqTgapdwPgLEzigqGreMowKK+4nSu1ugSdV8pvgFnJGj2BD7ewpJ8Z/7ViJtiFSk0joeRf8ETnNCnIrPgbmwwX9PA1Nsb5xw5NgH2Ec0qLTCmdyncY1n/CwiS1BBontniOHtXUbS/B9BTgMvHHJ72X52LvognNFK9RZQWt8QLb/wMxCGZG4DzYTAjOeKnvQUtb6VOSGJ4zHT69hk1vSNjYH7WUjrhown/QSl3SNONlkcHkjyyLr8RNdurKO+7b3TfbpQHJAxDv9MMDYjkQ6AAewoBrvXNfc/BiebH/UpdoxzK4OXXu0t9xbBojkFZ8nSBFlj2SDWYe/jcdruOVQsip9aNuzmTcA4npAPZl5BQ4rdmKEc0pyPi2Du1maly0VzOdYYn3ihgDO3vyhoVCRYTyEBnbr4mQy+28kH2BnRS324k3Gmmjzag6dcwnNg9Mv0ur04X09AnjY9cwAtTF8Bl/fSAYkJWDTO3REa/T04RMkFCcLMcak23wXCgvgmcRDOEjlFcOh9hMEgYgoV8Quk2WRAqNFnZDBV2CZFAVObwV+cd5KWPJMMFfuIhp5tdY6pre0vhRbW6ik5Bvx2NagEfq+612abd2svOFORNGoBQgG0BltoUWQxLqUbHj00bH8JzL5"
`endif
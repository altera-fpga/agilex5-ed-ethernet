//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Lg3VKZzETZrWhR4/f8SJexCBirdID5l+DMYEwNPTMxPvWj9HjrXjP5PTzSxy
KE26qvB6wvy6trIh9U79gSTqLzQuJNYppB95ydb07kdmoOlJC1KWcC9wBpjf
E9ikx6y2AYurZ0Fub6r/ftHidEYq5aotXksVGB37Mrq6em6aRJstCwWZ0ieC
NVIixTQk5kRK8yCuLx5qM9lGiowKrJ4yAgQJIyTVDs/ZmsEDUTQK2oFZHBr5
2hOyAYO2Gk1mAtgfY4yMCuN1Z05KkOcMZbMizwnCeYFi2FmhwI0S47yJ7XZS
2fuyrWUbF54o8V0IEH7W0BKhoAZ7sad8qsRCUn5Y7g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W5VOWxit9QIzpaXGcsJxe7K1k8VPSf77OcWLV4ODVYDVDS6O5O8O5amCKM36
jDYawyceretAuqYq8oaHX+GM5Gsdns/Tzn2PrXJ3QvxYFpr+4apHCHul85CC
I4eLP8ssD3H3x7ELMI20ooT9NdH9kEpIJU/LZz0zH/83TM2ZA6uiceoh3vON
URx6iPaBLrEffyZa2ubUvZ5eygDue1klJaWSp19s3esOHDVkvD70YMwhh0e2
5OMa3ZwbOQ6/s1BlDpG+YATgGrZYR1YQo72rNI6Hm9LJo7Td6dJ3aFKwzCd0
9xqEYdVg6jLAb3fE9gEazJE67NXPhcrIvbAa5I9pxA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mpF8nqr7sqBaGJoXvsIVeFRVgZhNTMk+Cz4N/99U9Y7oQPNut03ulFkpZvlT
KeKadLg9oruyMtBYWlNQB+Kfk/LssMGaLH/5ZGoZci/9nWCIAVr2ZwPT0FU8
Gmr3pPKMv3oRRzRBleF2K/bIYrL277bNSIYfS0srG06eapSgHnz3RUNPoHIw
qLK+3zwHjTgxdJwZf2imdjsfg4/+hNYRwAKbNRKj9ncJ7O7xt0x4bEsZthCZ
RDCk9JVZsHLFx6y0lJ0Atn5OPdOZIJEwXsMWbqpnSyVi9XXoOw70OevqkrnX
MS14Ye7hLQQeHPMtn0DExBxD+EZ/LZRwMfMpXAm7Dw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EfyU5qUwJXUsMEUyv1PYf7HB1orjtqECK0/PDQpQdxXCjEUX6yImzbKCh0cd
slrHXgmmizjC6LRx+03q479cmi9CZ2wh7/p6lgTUV1820R5p+PxluKbwJHsx
i8p/Cstos1G2F13FfKkGc5TtoKJebRHG6CVGhAU6nrEoFU8o3IoMeDc4/Dbq
cyO9wtWDsvPVkqIAEN8bi+FYrHi5G0iyi/MzU4GIwj+uB4FT2sF/FKc1CkGa
1oAWsACiL96YoZohbtq7mvt+diLwJv+bCi359ozFx9lTDyydJ+iirHsuyNAh
i/fAwysgDvPj5nfmgRK5BxVPci4A1KDkQiQAO4hIyQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EKKWNIxxJ8qrA2X/OLVZjPxmjcRbP9YLcGqDxTtX0IjLnHqlmxAAcdmZMeX3
pEmPHTfbtdwWzy9lsWCh0ubqLHgkkcZO+DkkH5FoFWXHZVUnII9ltMGnZhGJ
s1fiDOXYQ9zzX32wWxT6uGgpmkrj50LZx60UpsG2/oG5NWvaAm8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MrreHNQ9asg/NBgTZa4DRJVGjbFsltpGJoVgdA89KjLOknatjZ9q3cRyM1mS
wwlV3lBJUPKRPqLO/M7nEFcxMeWMVzqwl0y1vSvM+HixPU76V3sAOnsBZLkE
WvdWl+98QnGAXtZmmjgtjACm7j8VJC9pwzmTEccF8TAZSKADDCdye5BJT5Gr
eo+g1X4wsfDedlK/5lVSJsZ9244IjFqIKWucdlLA+wavf0rsUxDzQS3rUdDB
1d9F8sKI5xfvMBVYlUwqoR++gLQ4dlYqQLkKZMD4ZpyI6eTdE+713RxsqflN
NNXBSlDN6mT+KiQ8VK4tT8aj6e7WT5TOxk39d1QpAEO3USVSskF2NJctgn3p
ipRNUj3zMCpWpIoqVKYLR13/oG8rMId8SDBquw3mNfFxv5U0hsBRq8wPXlQc
BM6UWUrEtk5ZF8VVV1UsGP841mq66MxcIyxoRmwuI8PI5hpYwC3TWBUyeH1E
tmCfqDXHKcWmU20CrcWuvdwgAAGAWnki


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VM3IBmSWrK9H9Czs2ytrPUF/xKMnTe11mVlyWpfAAXh3FTx+m9hZGjMYz+Kp
3jetoBL/6HOXxSPk8tBUjmyZN4nblT+ZqQsIWBmZthwOYRStG6/0KSS5mLba
5w11zbDo9wDWhUmyN7Kba8EjzqxdnfbkczZ5nCt1qR5gUMEtg5c=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oxaNq1pMvr2XVAqctOxhVfuOR7kwnoclFZK6+hH3njoq+5KMznbZIKqfXDnf
fy7zzO1RGh2I9RUbNsDp+PubysklSR+UhRFIWyo0uqbCExHNmp/LgJZ1ayFQ
9cjf/nCsMs15uwFMIEoBGIWyfIu46h7l8A2mP0dkIiF9d6y7USU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27040)
`pragma protect data_block
htBuqi38hl/l9GLRVP7DDWPCZj2COovS6xnYwGDBvb86qORSMOgF5VJ/3v2p
dgHByOBgfAJ060lwh8sBNNuqHmwhR3wbaak2eEoLt90UASJkV20swCFIoA47
UuTtw5V78y3CWo/YoSXXNUNoQAwnOV7aPZlg5pMfhzNDGwNW5JBn/X8c28p5
qOTMoIMTLVhVzmOhN2DslRgfiXxLrj25VWHXwI90rA6PHztH6dgEn5GXtZKI
P5UAynS2oiofN2jBHaiqgdggvFvwkSzZW/Vlj7Lebp9grPldxOel+2zfBVQK
rwaAKwdXAZU3AaIj1JRoiXJ75yvcYyThbDpQAzWTuJPrh0/sxp6e3mubM8oJ
t2NEWphq/28XAZ9Q/XEb5yXsC9Fxuak3WPA8t1WrvvNODNqGLF8NAfoewi5R
cLg9FenmI9xxIoUXNI1+8Ne9rfh2FXnFG8MwKktipa/eT4D2uqzaPBWR1ewA
9su9RCREn8fTNpksOLHHF+dID0lWyFihXNc3CAvSklLWhIESax71olpk7Pbp
18vOe1kiq35xzF9dDgPMPKdN3R1HS0KC4FvcqxstG3PGOtjRT2KYjt6X+atd
IuLp55xWOtMFVAHaBXQoLMVL6ICo0yuff4Y/dOraqIpuTwVBgHylH4whiKjB
5DstdMd1geibaYfEQi9XyH6zyIdBQnp54PynOBXP3u3xAVh9wC0rT3zyYCKl
HujcZRCTINAILX1GxOn6OdLpxBSpihWpdsCzYihj+FvXgjKT/t93uBBrYgSY
BOJC7x1yMnEAtRjs9ilGzONNLVzlpzVcD4EjvrHPZtgSd9rH3HY+HbllK0cM
8exjz3zMTjZW6meQ1bPz7UomyPrurY/sEGU6PD2nb44RMhNIJkhDirkIsIEt
ANSJmbphl+0CdwdPi5pk9BdgWst4Q6jEpDhS6huMc9ere5e/5+Iy/xtMO7ST
5+fye/e8TtnSR7CwudctBm7Mu0cVNC7neqyvqDHW12+xiAJCOLyhvZ21Q4r6
UpQ+LUU6zD0JeKVCSrU8jsO6NgydgVl0KQSeX9/zeCp7QycpaoMN5hUujS2M
LDsBz+Vu6/Ah4GyNEEtjMNo/CJVWgvwirtn5Qy+cSAHw+sKcGfaJU9204cs+
1Ek9hle+U+RnGTYyp0DMFT8dzSbauQ3FwFzK+egDsmuJBa+2V+AciN4I9D/A
2L9yaW+KKcJuQBYigvBYwVxJwhRRd+4paRm2UcbxWoc3N2UbFVG1uRJOe0bs
VS5gg0srAroJ81rO4/61C1styzbhpN7SAnG1tadrpZ7/umhsybJotBnHSPoe
mBf8+a1HmKP1a+HISVJeZlE/xeSfY2aoPufu3/+Yj6BfNG+pECcnpqpEkasv
fK6BorvwaoxSg0/ABZ0TRahYL4CjYid35H0L2Puz2a67l76eZftn1SWLb2Gh
ZkLeIJOJdRAhXyDDBgWvqj2xVDoFHfUVCvt3B38snDSeCRpDqR9gw/+GTS4C
wikesx6/B8AF8jB4T7hwmqwRB80NoP+delqXo7/Fj9kjW1QmqevWd/n6n8px
wXnw5IbH42zFDrkL6OocF31l7ukWj/lv+b75u9JtMeJ3R923F9Xm1E81obGa
o3xQjIDAUjwzRrigUh5bW+PlhPcUJWgF638K2yPEcFKXSejpqbVK1i/Ex+VT
Gs6Vc3/79iocs3fOw/CcYhtQLoJzGb5JIx1VSuQdAhhXk4Ch0zjUbAPnMsTC
v7bHBR4bOcLCF4y5zjBY9DF+Zy6m8HKNYnviKbwfUG0X7xU55BUSBOA65Iog
k2/gGq3JaoBvStt2bfwmuxpmtCM6c/kLymm7S2tHuoc8Zf2aZFn7zHTq4NAB
asszGQM3s25gj2AgZSGMAwyfFX8iPxixbWqbjHjtEQ2zSFIMgh2LC4yNIoPP
oiWACFI7wolz8uERRngluC93UalotN1URzTBRuFG8x7ByygHwFtX5rtAWPQt
QCy+NiMcw+rLNPFvTfhFSVbm0Y+8eJi5XM4UsmCGQcmbJrOkP3awAxrBlASF
YUcSr3B1sLSZbAQ54k4PwEXPuIMapVGbpAjcJtDT/JwmqN3wddopMLHrGYmy
EnMYYHKPHWa5C51WpaPUM+6DPduRjEhikKk5Ri/l2Wqj3GaWiKdjm57Xnf2a
D4DosupbkwP7hJUgGhiX2p4RAoN7tOlYkpgLYE8iGLkhrfLtBr2vG/dTCQ1q
1Uuk2OiCmjM7FGcjaQ7h61BBDdIA+XmM9O9Bb1htDsVlWV661k7dLoxLMGKW
5grUO8kmTJ/pHtuKm5qr4u6ZUlw4zWFHVeowo9jKGNHSQLu2tv4hVo57yu7V
pva1iyT5R8XiT161Dbf0bYt81s41xEhurfFCe70/faYpd2fEZZ6bk5qwiBnU
K7hP8jQMqbCCVyRwdGtgRAjYlRKHE9/SDceWKATdMJHzuyAsOUNVqC5fqqkE
/wGHera5ocvu6otizTLRoSzFcP2xt/olnf1ysoSgnCa32IMUREK0yhyT6zC7
mQIU5jAek996EjfuMrO+c43LZTxpd2VgAs4ydBl+He6vLXU49HkZUfspIjKX
DBdi+Vmnh66OGa1xWuVtH6LNWJQPnNwMO8RnaZ3P3gJjHUiSnKajvBY8D7h8
iFKUZ5Y3AvnrCt9CPKwQMHGWPvNUc8fGIQmTMqIDhrXRGwmH9AK/PFZkxTRd
8g30Is0NFaKtnHEePZmCQ1WfAeeVhujSJH+eAt6CHWLFysX+rsrzpvYi7O/d
Dbet+HiS1VTXvScTUPo21NccJ+l6z/IY7n/GUA8tDufbwIonorvGpBTN5jSC
o8Vdu2QHsBO1te4K5HILxE+2nX4nOEMsSD/jlx501QLVx6IxNVmjVgsDmotC
c3i6sOSiP0bk2YMi5A82IyuTdcT/vTylmp/cb8JjLhq0Vzj9n3p7TMTWsSHZ
zZPMlJfgPayKHvMuFcTqH1D69wWMmbvIKykEWWxudEczl3mSHaOdGVRbucgK
nopU1oQBh33EV2ixoDkE3MJItYYJPPQoxT2ir/jbLCvEAs+m2THv6R+1sw/7
nt2Q+BIuwTogRI/mEZwpFAtyDCBuoTV3LGQZlaLPzAh1ic2EmiDwwinXCMwV
o1MzY2l56cq9VUaUG6VZzsWJLXAnQlUFphpO1maWDjgxoYPEheDlhbeweYh6
Evjh3MOyNYiMiGVmDIUyck6+ika8p+2iupPFbwh8n16ecJs3wbOR2R42KcJx
22y3gi65wNQkaENbdLc40ryjvKhqgF6pC/dePSdg57DelJaz4JhfW6DBn5Hh
kBFKzFcllqw13fYQCELPAd3MQbkj11hqpFPakQTgeAeJChuGUkNkSDpGtbnF
8FppIO20oyNnyTx67NNJTABXwn2vWYvP5i5JjnhIJ7Pfq4CA5xlvnQqjMmb5
WrxEqcOJnNlJjrzWRHxUsTg3N8bs9pHT/pb8v0dzZwUDuZUOPLC0p0DZk6TY
fNOkF3OJ+S4pW9IWjTImW9UIDALNM6JXl3zxnyQHrA0eNe06edrTSFB6taqj
k9gJoAWaAKRRg75q0VjyPICTFog/GLIEjhcoOh0toYNabx7CJjXMPHbjqIJU
5324rpKJjd/bU0twVSe7e/87CywJ/hBkugBbJ5S1FUGdnIZ3MskyeURdn6OX
PObaSvZdxWcpdUuZh1tGrvBF2Pta/V4min4vHoDplBQRs/ySOajr0ehjHS5W
hfCzsy8fLiW9r1/7k++h0vbDDv8tHCyLp5rWFDGuaNWcLO6HtZK45YteKBkV
PMRhzOaJrgUaR0DxmmhGsvCbTrSTuNVAHGaYPV7RKv5hNustoxn2suUwVjdi
Ej0KfegbrnSmamqg9++n7ulKp8l9GCkZD4VmTJh5hsjS86CR14BXS+49QeRy
HMw6DUSlTNguXAzhrR0nmMLDsxUo3zm7OKp9591mBQQUc1pqddy3x54aYjGG
i0VifDlqk0dtNMVfZ4wAcrv/Zb9jEH69lXcstcuRORuxv+075B7tlPPYm4lb
3zX27NUynqaqK5UFsjuoLCx8ZRMudMulZE8xwOcVdWMfkUEbKHbx7dGZha0o
xe6HVZL+6Xfjf9CZkpU4XNG4l5+QhbsnvcvnHyYK/IPqVq3exAuUzo/DLmvW
1CmiV611cvvH4Ds+YfpPf5Dz2DZCuqKWAG7QlR6Rgla+0b5YsZhHqnbR9WYR
boL8M0xgmhJ/bukDBo8JKJ8d+pv+46m0lYhW53NjuhZfEw1FmMuwLzcVu29Y
bbv3RoKg8UdflpnwnW8jpgs9CwQlkf+bMaRkhsUaEeUQhc3fVfSKTseGqhMC
qllB+dx+tsIVk9s3AYzPExdIrC4T4DC3ExVr6OrGyyIA8LXQrjVZKjAfhBPH
SW931Q4d/9JsNolPNqNKkZw6bH/+In54oTjLHSKftjTNbIM68FdeDlo1kFQO
gmuJG5uCMOsnFJLFFziKlFvbc7K0VPE/leNfCqKghBfYelRAlgSNtzZ66fBs
5xZrvIij8YstOK/7Ng/yYjgi8LwMK6Ob9Q3c9ge4gYvAQaei/O6z+9hq3pad
CSm6DZT0mvmjA+fAXG6n3UH2CIi2+GPVf19YLWGM5iyr5bTZ1/JptQvkdffK
TXS4Ez/3NByG5MgebpZW/kTl7hDCBGDCRgFVcpXKsR3NF6fCi/2yL2GVmX6c
0dWcq05f32XSaMq44ABWAFgO3j7cgSvDIQBO2fZBE0Mp6eJkDzH54L4TQcnp
AJhc0VNtx9z4QVTKV9sMqQLs3Ed41FatUly1wEUb/fFoA8l4yQh9p3nn8Ggu
LDZ7uTdObePy20DPLKi6k+hQOwMQNe89Rncvlmqs8DJWDh3zupmI5z/aURzY
M5yuHwW5gOMGScHGamHGUpTZerpKuXZK3saaU0fGlruWsReFYsxCU+2nchgg
xoKuVz5r66qtxQfDaRausIvuJtzsaF/4l5FP7mwX3AcHYefafml1yfIAD2xg
ERmNVu2xbAHzqC3jPGk/kY3XJyFf97DN6WCj7BpnOVDwrUAVX3BflTujGufS
vBm71ezAu33APZls6TRRVL2SHoJExFYtpeH3+RwTUPF1FLbGGMUIcC7Yey1X
6qJiQIZy8aup1HbrGs4qIon7xOJJyljq5GpcmGhwWkPz3klwTZQgiUBHDtLU
PgJuq5fMx90jpN1TwmRHywznleE8VCplCXxIE0sAf9ubace/i6TueDmSuaVJ
1RHdDZylEd0OkbCR2luC0XLoSrLybv613D15Tr+Gip4uP+plu+CpgGTT6w2z
fqL6xD7P4XB7d5/S6f1MMYzeEEJ7rWAzB8GJF0nyz0w69FFhAzVWwddxc0oc
pj5kag6Rg4j7CtsDpKsMgQyOrQWZzGjhUKqGQZBXFTmHVlIX8N1gt/uWxY+1
XADqYM3inwuhGxWfCJOAfFgLs8cB3NKzBy8Mj9smd6z4A6KPMrlnsdGjp3T8
QGZBZqAyoUSiYR4OiYGjdg++t1/q1I3GIYx8HGwdoQkd8dC+L0gGFjtc6d0p
SG0QTVNw4RJMBap0neGXw4ktMOHvk4ChYxqPN+CPv2sNGZ/1Q9GXRQCgmR1u
xsXE8Gn/mJbT661NZK7aw0lLxlx7Ql4eSybSG52oz6nZKNJu98W+T4xg5rqi
NbOtUAA7DdbBcMbPJ5LoL1NpeolCgUboHEmJBNI2uLovd6+4QeK+0mF9TkKD
duFvCuU3kaayYvgmtkI8uinv/kTrVlDDaQD5+jgjd21GW/4AY8ZR7Ig2V181
3e27Eixon2kGaStZwH5N/iRbq1fsEfIv9yf2tUDG/aIdEH0wjmLfV1SCmknn
jzaohMcUVy6qLPbXHpDOCrrxo1vcy6Zzbl7mPwqBb7hMKaqLCfkLws8efRAZ
oW0C14udJJUtNqCcNxmDVmm3thNjyHNS//7h+wBxAPnZiV0+P3DMHeKTNcMZ
XXSI/0hE0N6wm8IYwQGsmDK8+Mqb2eYtpt9UUKASLLlOlHO5rGYjgu/U0Mgi
088So1fuvQ7lcGdthr7ovwnVZP+dPvmTsbkYhr/xwNeElGIDyC6/QE4Zx5DR
faguFn51YQZI6LIvbTKyWSSjshFT3l55/hHiPM451E3XrOlCBRIoFIP8bhhC
/TLCp58LFgp/eT+9LTL3BVkybM07jl9lMCW1jjqsKoIPA025EPhBgu0c9jvc
NTnvggMsr12tofDoha+65wNWRbW+jJnrdl67DboJ2uUX7+TNx8i/LX0guDkp
EYxr7vmtkOXSNb++UIDWAoeoSFQqYPJHXsCMOfkueYeOWKDbYzqN5fDMXrgS
tiOEFiG8v1Ji+gpECV+MA+oLpl3VU3fqvPahLNtDIksjRUEPkvJx3Rlz1EZU
Ty3gtKMAptz8A8uOZWVqkfAXmim4lrgrHFPZRlD10JJL78dgJjUeBTUjTrLh
wI3ibxJp0TLZOCGsNxThqzNRrdUq/8DOrqKQUgJGUw1Ad+OiiJ32JGyRLMDq
Et465+BYRROI+xHzSOxDqve0lrdMyc4ch42jLv6QXPH4j6mRYbIx8K2ySK1r
kh6w+3SVfItEhS/d7akSFK3dbLrhXBwAEwgMTTrQrpuUsCBES5PtqEK/nkM1
gmhFAo64O3UB/Tnkkxh6ZlsO6ep6+OSDJV1e3P3rjNc6brU53gv2Z//wA342
Qsh1/zWYURpwjLqZ4Euk+z3BVI14csVLLbFU7gyudDoWskaxqeAq0oJpNR2n
g1PGS6UXoytg7iT5vGBnd++/+PHrMimmHlPG+zouLYgGliC00j4/gqrAecLC
ymk4k2WnW8R0OjNNdXwsQaW2MjJqN40baIvdhIDHsXasCBYEL3KJRKjFqHKC
vNXgvtrJA/7qc4+0eInf/pr4N84NE4mz3bwT4Z3Hz7v3G0olInJlAyDYhvn7
4ESOkxD5J8N5yqNj8mWfBxO4dmpue1osMAVyCTVY3Ryf3Bwqj3+AwXY3Qe4Q
o4Q4X2p4+cgkakUOe0Dy5tk7Kg612DFFYDC7nt5yHVbbHGfzEe+MNju8ZDyU
PGpS3Dl+LQGKzNQDmbkjDYsxDbRi7UhMQisEEA+SdAk5b3vWuggLzGp7hXB7
oN1hUzpr+Oog0QU9sFNQTJ3ew294b7ed6sSi7Bn4w8ozqm7kRA3byl0GBZsd
LWfkn3qdWOYaHnvS7URovPDy+ttGNd5gDmfexLgGm77EDwhk6b4LTrQy//Qr
DK6rGH497kzWr3/7b/Ke4CY61iW99jwDo870Eg8gEsZcoVWS3bQ3LxbiaaU3
Nt23e8y+C7F76nhgFzp1lWfvVjxOWP9QZfILMmIzpsg6DhF7YOrt6DCmULR/
wEVAiqYIo5ucmIFNGCTM6f5YRpPBnf7lST5/DvR2vLwjDewUm4BQ9hU9qPf/
7vxWBx+PL9Aep68o6Rn9E4w116mP4l0ppHHGZaJa7Nn1J/2pDO0Tc0zhHpdc
Rhl0ke4N/eSlK+ZOt7tdg3gZXJAYdmnThQt5SstUqx75G8O8VNeUycH4J5an
jO0epfWJpfFi9LgnUnBv1R91Lykewav3AnDCHM88F6vCIPF+3HDlgmQA18Ao
/RPBWVRMtVqWPLqTEOHx+CExjWLtYdbPM+S7jGriMC6zfkLWsyL3Z4MsGtyr
9cOWU+Ytj7e8Zl1CxJbXMXSJvk1gS7qxwrrwXONRPPm9qLgzo/f5wJmTAGTc
Kt7g+QrJ0ROCqGlQOWWJ+H44hbsCvU28GU9orRvfNQwPBBgLB3/I4wbYRDzg
5fHv4YpIzgErHSOID9JfMKe7GtYEAYvgVJhYDcjU6uGI5HDdR58M/SKY7QXJ
QiCZJrVroLSAIRYeCRGvqlS5GpVitOkoJCHtaUK0ser2vyniqIveMY119MgU
9KaJopOQH+qO+rezTsgRptHHYDzZ2E/OX/TLjisVnSOtEW7Pmzt52++aQoZD
MCK63gG8gd5BveSR0LS7D/8uiDmZZ0gurKescKOeWfIBIEJ+aPvLMuH3Jx3j
cuXQNF+E0RqnYEs8HIpmmIox9YrDCaPGj86C9p3rKiCGR9mIi+vH/5cyNvuL
AqmO78oi7PNALJtBa20+huIuq96n+GLWtskoNp2vg7fhEDa8ilgg3R7y2a1T
W9QZqSYydC9TjqRvcLRLVYiS4XsQkNNxwyrGSBH5kvBjs2xIdYGYJCMLkGD6
lIsYC9oUh2LclIJI9qxZ98tpwcc7JSt9Z28VKpG5TNOa/wnbcKzi72K8KMY6
DX4kwExgbqLLOa99S9HKOfb2Mgi1kL5CX7md+pOyAHqJaRNWCIbiTMyrx0Bj
CNz4yFh5okItobMs827bClEeJ9FjRkjWGNf6dQZJkyLU3c4oF6V93GNZlB7/
9t4chcJR6aRK9nKS8SGR78TiwpOQ4OH8UTRbGwHJZwcO2UZlmUOCazV1KHVm
nFuzcVehfqK4ykWql9TD4ZVtWXACjOuKTGz28VbggitppyvstZlTQU/UhQPJ
akQ79F1x5kJosh85MJ0riA4xa3tu01MH63AQbgwUkcv1iqEqEXn1RAUb928c
6SlkkBjZnMfvKZY6U6V8HeyKSjMYJCulykC/3E1MZrLmDmCbk8KYAUUsVKAw
SMMWzfgrvnwZyUfbVRxrfpFQEU1Xoci17n1fvt+GVoWa2pieRI8sqPwAEHFf
8l8d2rbFUl3LTF4GMnUhz9P96TI6nQrJ50X8w+2UqYZaKrfzDWU8/3SP0lnL
KsJV5HDboCUJYEIFXXyjPDApcaoJomx7UWKTXnvWbvjG3BK4EC9gpvATQQkl
kOCfgZ6GgMmM/cxBAFaKIYHa0KAdIIzRUvg3ZOUHd0jAYL/xJoOEWAfxlwM2
CDCzH6qmn76A1S8+fnxubLS2Q7ByXnAJWf71rTlvj+XzKgirvGE9s1cEVAMX
7bXm3D9ppm7L+BMbwhw8L3zCPAUroIbVQUEGF1tvhHg/jTC0QKQMrP2K4KrK
liYgGWyH0O0a6iW6H03DsjPWaBjS/frEgmCmeHfqkKNe0vsiw1tAPcjNP43V
1iDTh6pl8vYemZihAgcQ+LnHYHZd43C2xBjr+YB/ke3INb4xtG1VdBPukx3e
Kg+ZrCkc+FWdItsZnneRXfiADrCwME1pxt6LizYrpoZCqceO86YhvofqGO1G
oi0wU+1suv4I1L/yVRX0sVbrpORrFG6MAGJPV0+5LeGbwnl4K5wKZXr1HXPg
Y95TNN/ifTXyyGry/3Ab32HsNtRW1oSiMK+gH+l+9blW6BnEyHs+QayA0SM+
VBmboDu9sNLxrFtOk6uNSzLCB+cX+OWdcGVK0KvJOODjLVFU9ysqzqC6bI2A
Tq/w7yAGbOTXSkAzXgSw6tc9rdRJsAbjzx/rYn+5EOXuFgPbwMiTjqvmGEcV
zRZK0vAM9gZ45AvVdO9d0Fq7H4wmDbftws7kcBpR7DTnsiyGJpW2h0aiMPOZ
njMc0xVUGfG5B4n/bzL+W0MzLICFZQaLg+ZPOI1ssquQgDkwohrF6shCZ3cc
vRpDkJDgJ2JSlwo9bbEVlsvCf8Ck+8+vgcqrlhD1OlvwXYm2YZ3DWjt8UgoS
7SyKN16LCpvqqUuuQ6Cc0AKx3e08tmqQWA28C8wjjfjrXVt0YWyJQCy4Iyp+
1eW9WFU4pLSRMQCAUHJmdEfhYCVd9gKk4KmkJo6UYiAgSFHL5DSHNea8Bcyu
92yNO5FDj/qJS5mKmGxrIBzUfpyXGLUfY89chYv4UjhU/G5QEyVM37nfeE0q
5xe0s4stitibIDWLHoToywEvcjR2jOqCvA1u0zPP93Ma9KQrt07wjIyEu/ln
O1D2Vd17s+dNczdLVHh2hBwYD+9zw7yNTY8y5SeHeuUxkf3mKW7cLznyx1FO
tbQVlR8hDlMHp2/JD5uAppN6AmPjcpgZTKrPGwjAeRhTLz/mO1KSB6XHIJMD
+PPlEopUvWTPVu79Wyh08NxlQPEDA3Ba+urmcpqWNUrSlcbGHAbYu+7C3cGq
jMYs4hvGJRiJ7iOr6FIaRPOsZegSs5pbfYmM8CjnVOcFzuasAf9NywAtIIhd
lb4HapJmTmuG806H5UdzAafAFqkg7KjDCEaIZ1/McwRdLL3sMeW9eeNRXT1r
bdxaBNKDscwfpsHSyr39GQj0pmg/ZjIVY6unE7EdeFziT65h4Z+U0BpwS92F
4ocio4ZdrpG+YMUEKUVb06C/YzbaYt51xlRJW59Uz6KKqZHrqVXWORkCRz/Y
dr5MmNj1qqRaKF6nJ/OkcSgPWKnqSeSwn/6Mu8og9EmQtjkgwhMKS3RvIiyu
f8IBmlxSMLVZIkmeVwBqI1bVJKfFDpT/y3CHGxvEbC4oNWTX3584Yh2JIhPN
vI/hucsEb8yfPOOz2ZyjF1DVx9IZisEIIaJQMsc+ym9j1rw+NrXYBQqGpIVJ
GGrsHk0ymR8w539yLWle+sqR+1fevJVqL8Gw+7chXCoR27BeijojzmvSpIsG
CT9yDhHmbGyyDwVPAcpS5b7Zw4oDqG4TAsheve1TtejWeevRr4dmsysqizHP
o/Otx4b9KrWzum+r0WKWtTqGxcILGqsXFgf1S1zqV6M6Dk93kHjm+Lv5NqzA
QLsWdZUkHFnp+tNlwNsMJRgpUU62X3JyZXRchgRGJOyGOL1mbEmkNZ9ssFOK
GwFzk7vESFdwaaFRFQ/Gjx1mHZFuIC9i09SnIB57SXeU7WiT7VBc7Gb1vYFe
qb/6XSqR8dqSp9+uzlkxAfjRYL6ug0P7hdCOFhTbQWkxyxI9miN4E206iT2I
662XjzFQxQf2FxEpJo8R4shDcT2kHiw+2dDBhw9F3jGXUwhahm3aRjMaD6El
LTpHYill4w943FzPg1TNS2SUn4pZaFu66kbgRx4rljQekbHcblIKMz7IH1bm
ZsgbARcIvAE4gQrA/aPexGA9t65yX81Fn54sCmLVdXuElAGPnZ6ihNnTL6PL
TwZhVutEPBu6cvmFSctFTg9DQ1LqM7Mti5zTFGjmapmpDlc0UDEzNnpqhOM8
S23QaoGUgix9G4xGrsDQmIOFENelMh2ol78q1w8hSFQhnCe/2R8ryOhS2hXJ
CXx2lKLcmye3jts6VzZCxUGwEk6pdgdCGDsDJ8p7RSlmrHJrJW5Q9fAMiFWF
7SXJTdWG5sJODqEtG/PyyBb2Ai6JyZLxtFkm7fr/Gsz2ik5ixHrLpkm6bOOy
FrSgJmkSFbRbMIV71n9JpdkcqMivKuMlO3ueuFav+tOuUqpI+dTYeod0wRnP
VBRS0IEIcwYB4m5ctlnXNWk2Ioe0ehW3WBkelFqC3eHWbRfScdo4BdrQ0Fyp
6o7FPykhU9whrqz+Sj+EYpbv3Kf9TsFHdckwPe3RwEO9U1JjqVr6syXKBsF8
lXLAy2uG0qpxo/rKxxLm6HzsrgRYf2m4OuEGCLufjFXbww46Sviwp+O12OPr
SBP0RtW1MX9jDtuRXSeJEIfR938Rdh0o58czQZx+toZ5/RQs8uiHfdbI53w3
304ILLREBI+oZu+TdAwheXSLE3Js5gacRH/oG+OGesUJdQm0Cy37lzxQMCI+
4l80I9LdoCkjeVJfhY8BrrPvg8cKbjPA+gjyrQk8KWqIqr6upeMSt2egFL0u
ZbP/NMJL7K+5UexjVBj5VIkVY/wvFW26M0kPnu/9vKBdKHTbd/fdU/0HRqWA
POCI7KUwNIb1ftgKKPQ2UWElGoAtNCsLvoT5caljILOOTSeewk56Ci1uo3IM
rP70SjZGI4TrrtF6kZ85WE1OS9RQNT8l731IkfcSlVX9fsPJGR6POUIDlqee
9Kta1nsBVJOhh9dhocrg7LrxLFeuR/3YwiPV552jBAoRIVxYOUOaQPtDN4aP
sBh7oBG8eIumD1rG/TnxfFP14QiesuPIAtEn2fOvUcQt7dLXsT7S/hcvFcuU
4HKA8viKUzjWngdDNrJPso4MEXpLBcf4jBht8Lw+7wXjCXKZdgh5SVHzZIiI
K28xNlE15f5pnr81BHojG/zzeWcdi+HXT44RtXHNstlwK/Xe/q5trTevt+sf
d728bVMkhsi9geEP2hbN19uafs7ASNyukmCUHA808oy3qIazIwqvOdYKn4H4
ZEceLgic70pcSDBT767y5DRt+NREUXMDeUeu+k+PIIpnc83x1K8U8eXo+PR4
j7m+KwG15IRM+di5FMzAG6YBEpalffE66v22qG6LXRoWHo6pQ9HvOiUGTrM6
K9n0L6n9+0M3H0FbKmizc6cYGVuv+MtS9/qs0/1YexwuYlp/jyiaEVtmr9yr
SMnt6euCUmmYYrRUKnNESNpgYoNIucGN7jLLg/bARFf/ePnvSBTx7ZjgS1/t
rUBa+HgmYbSB4uAlO+wPn7u+7iruDyh84Jbnn1yuO0pYyGERfpFrym8Ix5Aq
3pnWCFM6jRVh5k6EheAtrlypvGmAW7KK6Qu+fOd0xEyxU3yra7Jw2JkrXWwk
BsWldrupwQ2+v8wtM81OhFLWQn6RKNc7oooD7Pwo/2BCYS7Y51xqN0Pkymxv
RbFojeTLT3KLH01IP9m/35VYctrcjrFU6eSMNaP1wMTyhvFZOky7nnpZO/iP
6/31aI1qIWX0tfDUbK5rIiQ70UVebmlhsgHaPwTCMCyot6weKktAcwqRRqgl
q0GPRJlCZ6Jcuj8TvoU61bf9MR1B2X3V/6chpFwJ5AymWnLd6qauykG0m+6x
oIldHi57QS+xjvctx7fhkIAVTWC/EDROMg3kGmTjGe4vQWov/GxXLwhtfXqG
kd/FgNUJsM32s/g1WF5GxpGTGfBT0x9x9MIPy3ud5dxMJTRDh14mjQToFKzD
iNEEKiIDaafIhW1Qkc+21lbzK3eL2Mts0tQay8eCvV6mFAfPwiQ2k3eanexf
Cyt1DhRGqNOvhD9sRxn0YCJXmjn9ANXKFzyUDvt8nJ5Euszygx06pHnSYZ4N
Qqrh8hB61TIiQ5Aaw6Ir2K9GuafZbcIcIYjheYCrbG4D21eJrPbnFQuLHViL
Bp7lT9tUezlIPvtff8jlgy3wSMSfIQm0Xn/aew3FllmznQe3LNkKDJ2m8tpl
AbXzIURCDyYhWYKy+YOH0Iw/3Ax9SHUVgQaA4PfrTco5zXbMzp8uAB1eb6fJ
9tHJrFDNfW7fz+CsNvI1LEL2cVkbfI0EO+oLOC9PMqeL1Ba8tdC8SEfziOYX
9r6GcY558E31Y9cX2wIbHpZGTYWWAQUsZoaT16DkAOMk32Q43Mu9Bj62xRwp
kDMv6mo6sXw01zzEeGoc+o8a30CHRzJOILJKE56aTT3teTQrEIYoa2d4hJNy
hdkjm1c7PfmxuDpiMhKU8b7Pnm9sB/HPV/UC/brcqa0BZltfHbwiK/7EdJC6
qxcaabTVfLEexiBgeZyuqQRwZYhNxax6Wk84z2KqNBOytzqI7xks1IrVPV7U
+mi4opOJeUejVYHFSgeRo07+r8Mw7DeGo1e8ZrFmU3/S/nVkKu0mX4msar8X
J0BacUyrkIDYFC6Gh9bKGUIRCaIUeR5DCgzkUTp9r3T7UiYc/1eg2i5VjD8+
5HvlNYKae+sThTXtd8fo0Kqt9mO0aVtd01rkd2jj7x79XoOW3KEmWAZn18DC
UUQx4bFcknyq9urFyebZ41PpNWtqnvw+n0bZM0lfbudFwTdNUjxJtmt2/oGt
O93XvXBXA1OUPYG96Z/Rmjhq7PH3PNxDjm3bALpP9ssg+yorI5K1j364+dR6
rtOmDJ1GQ5Na9mTT2R6YHW1G1XdJJh8tT95qKb9FUesrM5RCWeVvTvDwH4dd
XDLFW8fbXDY2fRfRLnxU4gCZlTqiFaFo6+60L83Vu5gc+WSA1WuGDPoWh0qJ
aRAteFoQRX71zFow5usziQcpaCWGxtwUsUWLWtVKb1pW2DbKVc613RVWKwvF
nJFBFYBYNxF7uoOJJ5zlCtKjUiJ0QkzfOi/IqOA5mqeWoF40pyjfsPHllZn8
hCgvQY4JsLsxT5pcrEgt9j0eEAmxhZbneLXHNfk1N9zT4vaQMShGjsmYAX5k
YIHB/W7j/4SfpNIpKbnd8eCJ+RaKPs6ud0o8daxMZjTji3kowlNrCyYdh1T9
UHdzeEghmtetGVdH/YHsOgursxqok03Poc+RTtIOJhEhRU9Td76ehLA/3MAq
ePn53+zEO3QwJzVT5UEgFU+Km/VCg3nOoR+84UsvEAafVT48Q73AY9NXRdxB
j3PuSUO7JpoHaMFSs9nS/gDeESyiKTq9k0kghUWnIirDYaOtMNjriTNT6kD+
7d5pI7QQcffd3W7cXHZTHmnmv3Z1kAiJDwwR1sXtQZ/cT36g1vAuasGPevsu
auHToat8Y/kRfzTLOFkuZUxtqrGKNfwLLZ7jsHVSWrNX2edAM3F6/yAi7d8W
/vlcXqQZ+xbRNEAgd/oHmxDeF19CKgFVhmDraSkRiKaRodUKlY/ewvAMtgLK
YVOOOJiyGPnUgFoQLAo0VcZVQveWiwCmCihh7dwKGPBRgqgDQUEUhqWHzcqS
8+ZxJYMfHE+zsqI8pzRrdylHdai/KgzU4pxKF0KJ+6e5d+1DRvygyKXIwsus
rBsq6hC9CfNmGfGiSR5ICTcpR80P+xhVeMnoKH6NmwLRpXAmoASz9lc+2hM4
YvB+ciee1D3trmAjbiLDtTz1B1saPj+QgSHYzSPIZvNUYy3DaAL8U98pbh0K
0uM7+w92Qs9XqFKkxZynfhtM+ACIQH1amtsrdlNiuHqbjtFBrJZ6BB+wtSqw
9Xotj3tcfiQb/LjL3gaBlsL2vjoEMhFVG2aI8bQCA5YOF6QxYS02CRUc1ywk
wqOM3NSQiACqr0Hema+gdgUmMTNSc2EvYs2dRT0wsj2iokIABglW4543xsGO
5rirwoZuyHvgAbEDJqB1TcFSbmFhxnl7Lh+qZ4S+4rfHqWiXEz0b2mRtcwn4
5j/34CgjelwmKRDPtF95AYTGrc/XqtpglYErxhnhpsZcrtxwsbUTe9HrEEk3
hljUFor86cfl2PFKQnZGTNkR4MMq/QpGNJdmJb0ex0ADvUuJS0qkVdi8Ub/5
yVi91wzr7RsC842bs0i0yzW6p4uJFwmQ1zH3waOSZL/2/DGdZCqtNfQevi6x
TLBjGa1ahCYA9D9nM+dqpacvJcegGAR0jFD5kaGakO6PBe3Uy/JItsnPI0SW
P23jh+UYobmAJ9B8W/VPZMmB7RVw2dTEbeWVkWmjAiqnguaskYned5HylOZx
upHOQ1gO/vaO5q1VHCcSurcg4OMyHSyOmoo9LZQpYQSh6yv5WS6lvZz90m8i
A2jRWz2XHVG8ruRGLQTcOdsDvZz+oCqk6ovsvmXmquRVYzk8uI8MD61oFeFf
5LducjpzezM0hAu17+3hq40MfgYIh75YGaXSt8U3IfP/h/A0+VPKetADUHHy
ZID+Vd9LyXO1eIYP5mxzfhN56d5v6WhxeSWjrAWwvujF2IHJXVMu3fEBcZNJ
hDcGU1RKzYDxHP5zy60B2KwbIbgsrjo37WOzyCbdZ935L4pF0RxCabLzrdFD
DIs67pystEvetyyTfjhf5bugrt9rmVh3M1t65ws8m3XI2+ZVi1GSRMCRC9f4
V+WuHXqM5Kth/HJej8SDZwxfGXLOTMyw6AlUYEpW8sda1HMZyKqM2hslex//
ADsB1G9rpNOtDMSV7oMH9G6eWtRnGSbguu/HRt7jEvkcGYVBjqWnIWYESGQj
eSNzKuT3ofatrXly7qIP3W2wFtW6Apn7oFrSz3t4VlfoQImwrqoJ67uQGqT4
YIfz5CGMteeWjvG7GjGz+XpNhMVNYhaBAAevezaxByPo0WaaHOC+knDBIhkQ
ghoFs249e72xCUciadzMGj4MQVX6U0eWayAvaKbXtnYBMQtYhtEO2hMA1L5J
JQZz9YbHWDvOuADDyRfQCRX2eWSVEOgsUs/zv672EQYGgc18YzjaNULl/CQ0
Mk+9UkOBqMmZx+GnNzy2a4sm8tG18C8OjpiIZBw48DiJl9LnQw4ofHnC2FlI
jWRVjd+0+T6LTDqWpkiSHsGjMW3wppLZgCsGqm1GbtyHPGvjepk3t7zlHPyP
SlIpNWnLunBEGtFf2/0dlp4awUb1XwAtmXZSdFjE1KqLccOg5wNKAH2R9ddp
NI2dTiH6AdNmDWxeG4T0LzEIa7CHJ5BmA18N55Z2PNpiFz43bZ9gsnvirF6Y
zNU+uixKS/Sq7s/+gsKLktdwOrNFV+7NhHG7flykEKLpRQ2wwGKdvPt/XH36
g3Kn+727dYZEUkmc+2KO7bRKEat4cPEK/EpLa6NEeaQGsWAEMQuM3KIayOwq
elNs+i/pT1Hhs2goqAdZMmv86my5pvhME+6C/Y56RsysM0gKf6N3BoYLNnJI
z/qHkd43ueIBmJcJVN8m6nW2sqR4rSAiiiXwfYKWAYJtiDeKGh9Pmv3gIMMA
/EYnx636qHlIQK5n6VIXHkLgWv4z9Jo4yrIQuO1KHhgraFh3pDt+COszUFzn
fhhGb17jM9rIRxSmHUgBqLkgfl2sL86BRUeTvGWg59DBU7lG5QeAeNwJU4mb
b/HvJfhfGQEDY+LURAK/mhNMA5+kjz1otZmc/Vu+tlTE23Gx9cg99xQtRLfx
65o/xf8rKtnoOb4EwSOZ2KcqpT/ZVnfBASByslHri2Xxgz6uBEKJpBLf0b5c
eEvogml3BMWXxcC/k0GS6jjW8kmTFtrWW9qKte2gE25jTRTwQ9/5BkJLcLUt
MP15gQJSQxQ8FPYHDeXMW4+8LWf9RG+/lL6UZFgqH9V++f2SOH+4VT9yyWKk
yTaLUSyT6eefYerXd1GpcGb68hfqNZP2DOARzvrZxELWFc+Ju5t31lAlX9KB
ftNNvQYRmu32XPldBZaa8s6j8yVZikZJZY36Z9MjRbEvhxCsyFPQhc/+ey53
ZJAS5/gC4EX4auFSTLp7n20fhhzN/LYqU98GlroWa+d8c1+BTw251QFHYrz0
X98Kpv3kpJJLtxV70fTMRIKdwIRytUmpXU4SHyFx1dEr2NcJGS6yQ6CpZrEQ
eYxoRMD0sVdOnAyEymgOzUe3QUd8dpieFyLpX9n6WbBOibY446AA2wLgO2sL
Ek7C40pDrmzstKy/HOjzw781HmPz/kIal0COK55hMejEGpmBDU5Eyer17XQg
f67hd/R97zlIDRJAgiOR/vHWsrmUoX9B6nG7mp8nlMCu+NF2qtsc8NVFy36B
P3Ad6eNGU96uHibh3sYC9F11bQRCRz6IpvtKW/DgHSdts5csQeT3ODIknnfD
+LTVCwekSNV6yGjsz7Pm4A+vrZZxTjao39OayzWSwKhPbd9JjTEvtwIliyc0
tn3JALkuzDmNnreb8MgMQp0snNzcDCZS0F0PqXOaueSfXuSwuArevNJNLeYl
NHtozWTjbvl6mx6CZhwminD3o9ejLtsqinWZmHUWC4Z/t/l7ma+Syqw3E4Cx
JpgjicOCwg/l5aeMhvv+bCL7AN3vsja+3DVQ0cMv93X3iH6vdnebEF/pHVh1
oH8GE4T//3TRUDSRjWcC9s5Jdh6W5SoqaRdfwU8acqKQUFFdC+HNy7rBbJ3x
JbNQ8XwA+O+W+Okpec4huDaJlrzkc1/LJDjfQ4i1dv4gIYvnk6/bkz2yokKg
IrMtaqeCMGPjg53GJ5dQe/oSNlmG3Y/eTvb6n1VEn+j6JIHfdJdBxTzthhee
YedzZ//5Baz9jI1GpGKsRSe2t9VuITSP24VQSsDgoYUhzm17wv98KEN7fron
77ZdjEcqBz/f8QpEc0AhYJt8lytYR0b4ywSsgbDYBtqXPJd+wjS2QBt5wEjj
Q10RmUe+0O33XTcMLpmdwVZIoBTM39ezcMEgu6HVnwtJxTG8f/CR1vbWRq6n
fbXxl+nZQwR72y+LzytOf7dLAXSvd68QShSJzCbCPRuKIGgKHkS0++qYZVEJ
eMohZLQhQfbOJ27Fd3aXXS3+Kp8QSKYZfNxU523rm+8Yvnm70oRah1PilK9v
/dQwh+9QqVmMYoWmOZu0He7ILTLtx1w6CEcMefgIIiClfo6LKL+px3I53AIM
DT5E6b5LIaEdTeV7/6Ol70IOmDG0uSzYliDEmpp1t/NuDHvk4qr80Hwsu+Y0
Nepq03EFjr2VRqoCbzaMEkoGUkBy4XKLFr/wSzIdAVDmrmj7LheJRSQR7MOE
Jyi3LxHMh0QYQ7aO0eAoB5yFQ+h0IThq7Nn7hPUnlmSeSYUI5BsNNazHI3D/
Vl+hWj72bhr9mNZWmK4tpQ7/n9/doPV3avMHOn284MqTVNcNkTO6+kAPvOpG
f+zxpmuBGbkSPZ9x5kVo6rR870BSz4GwS1BOYuDx+7zmv98qJMJvgLJ5NveW
bIKWUY47Cc+mQSSYiMXGAtVrCbbEsjTveYry2OePhVI2X0TqIitnEDAnXPfW
dEyi2+mhQZenoMIJbw26WsjtEer3XwSGYgORqqIhLqXzH0qacv2gLBT5bNY+
lC+baZw+G2inqjAvzSMQfGVne106vEOEf9zOrZKqeysdDQpHnw1kkyG5vHbb
A4JYe8dhUOWN8Hw9mOl/ir/9UZX8W/YDfmgIdVQCJ1EGeHipwdKV+6flZENd
pACbjfiMN2P5JcNobKhj7unl6ojrcBZPOgUQzVeEPRl39wjjQbp7z82hPcV7
vil8xcx+hglQXtyklH+JpT8GuoE81spsQ7eNATgj5L3mcXaeuyaaeWos0Skd
oa6NqDa2onvWWbu+phbDz3SGZXJa050M7RWZ7Qv+73P9SjzDjaGjSTMYtye0
7zLtfX3KCH+IiFggn+ch8xt1KsGp7ZPL65zcR0zcOgVK8nFkJE/YQD47IQqb
16YEYZunQyLN1d715hNDdD5j2o5gMN4yQqQESC8Qbh4zMS7djWu5/hk1LOvZ
gnOdenutmlqzuz0wZl5fBGknTaqwHGrrhTT8TcMHsKFk1Ax2dOlFwg0w2jqp
NdieSlCTFPGScidWDcP/NmqBDBW2Nbs4a9gyVf+4+DZTBhBRbLnVCLaYLGg6
/lP3k3qXxGAOS+JKW3I/VKqAK3D7cosfw+CmG7Ukp6wEhLeW+ius3Iw5wKSW
YFxSpeQlW6Om1zrNcPfPxhOEpxV4f2Il//j/m3ADunnB14DlSpE0jRSSXHFA
TrPJJa8qdPlr0ldHTLMzv0HM3gZ2FbiWoE2+4ooBsXHnuhMmyotIL1DZs2Uo
yq6kbs8jEH69+bJibGREr84N8arv7yMrVmI4mZglKHL31rsjNqDDQxlQTeY7
DnOUX3kjVrtxLwiJFpKbzLIUDBjaixVYwN53pDIWBPAthUSSx0v4mNVO4sdN
8jz/UxbSophxbjn3gG59W7KZ9Pdj8anna11QikT6tBTQGvV5DCZlICtZyP+2
etzIPwxY2J2cWsoAvO/UR3XeHGvWgPHKof69KVcXykizcKZdvJspZ4Fkcp+o
ghWs6grdmVCtSFthgu4uu//dHas4r/gTc52amIKXzjuzNbGXZm92QtT8cZ9/
fz5/7W6Qcg766YqSebyVMbJ7OV6gtWU1MjbaHTlNgARR5Mj+3R35IIzOAOwJ
up0OXN2Denm48l/21+Ca948Vu9Y0fPrGkjybFIybRdKEd5IgsylpSRmSOWOZ
RK2CKFjo21bhT2wVbenz5TdEHIj9fQFiLRoOILY1ivuqqWJ34jZ4WezuLPTs
35VVIQryghh/VcuGPJja5dHrhWRoNM1K4nBUJlseLuBUm8OQz4aYDb2CnyDB
6et3myNsLOCu0nHd3jh/OrdUxRShyVwnzydpKy8S+RPTtZ1tlcOyo/P+Ps4Z
6BioLNx4Ax5f7O1WXkXyuRQwRIiX+jwCBrdYbGEl3Es8+9cC8R/BVYtaYjm+
DPiLR2h7ve89YntYCJupY6zHC1JXuLJ1zhTWT3DujAE3dYFh1JBaEqvMKehY
coG89Cs8FMTjG0JlMM3pcpnADc4IGRA22lTAyny9lpJS1bLLonu2rgzqWqAm
0AvMhDdVmHtLCdpbeElfxw4D7PUBurhr9nhB8KC1LrYfo26p3r5t/pfKWYZq
COn3WKF8CYVmHogJGBlAycVwIvWNmSd+ipWenLzFCUmWI6TeFvRVTG4quQz7
Jy7HQ7pWyQ8JmJ0XACgtZkFDFCjdvI211QhImGocwovA4ZYOX9c2Ynw9syvh
YpcsotwfnGNEN8m7aHWItdv8DM1ARsMtL1zcCYf2Vh2jj5H3Jb8msR6it+0k
Zq1DvEU2v53RJlZDTghJiq3AGQ0Bm/Vaqix/sx2MwL7g6AK7PonSkFi/WwB5
fKQsgkD3c4vOZf4buGeHmusP4xO+5FJiLjvWPsu+4MET6XQ2nIc6MEydt1OV
OYzwEg9gbqVbWJVcPQvf0Z5EKFa7nqmz+R2bKOjrCby+WCveRIwfqcqrVKX2
jo0T9FVcF9NjDMnkIFzvy3y3BfyeVs3skxLmoIwfY84mUy7Ajn9PlB71EE8h
L/5ZKVj3hX52OyhjRVd28K6f3QQ26uRvSnKlps3+reJaHYdj17LMLzzET7T5
y8wHsBAWRbHzW916G6NOPCt6IYZGE3dWQDp6OIF+C2EDISo1iuDOnFgKhOOt
TXqM/dCiKDS5aSbr/NnZCShsKzhNiUmHPt/j7eLJqoU9ylntHRAhEOXAc/XE
ffPT3kpyoCmfeGUxpMfNvrOe8OYlmbPQirv9ap0XqyxotGThcZ2ynOCYo9fv
7XwkpYl+I0ig9hklFNvyl4dJByBx37BvBW0QsHkcEoEsBu87lJ/Rz8Q+b5WD
bb3xxX3kVsJrpBY2WFJMQ2BrctHL9L8BqvVudV5PWSwwIwLGQ98uNIoGtXv9
9vdtyhdC8FXk9SxFpDFUNCzVEV0W/Pa0zA0cTN2oqZUefUFrbhu5MDT6XwQB
ujHHCKITY3vXH57DOKiT5TwnLKxkrZahFDKdE8+FbJTBA60m3fZCnsN5pdZ0
PvtpCy3+MxLc5kDhhzl1ydmEoeZ/61fdJfS9yfyghieCmWzhDatVOQyEjqUh
TcOsldKZQEHnmtfm9roi8/y7vo9p9XkpbdWKVRxec2dq+dSwHMyHUUj4H+0j
c5ZUry/kexMILNL05wrYe1Vt9I8ML0JoGaCV/I5sHMBZuDbPB9M8PGz+nadY
SGro8lAzqRkSlnVoPNXU6WPv+dMeJLZ1HNujrGF2+uCKDSPQRdLfnBeCpyjS
kFrAK2OtR89C+x7kITzo1VBDH7+UOCLNBBLIk2LV6TypuWJeMf9Tj8T01cOJ
Dig9i119e/4ios++YNynw8WyTY1yI5NcfPZPLgnqpGdpCSOxTX3P7XPENycD
9xg3rMVwKn+r3E5KC5in9+9K0LqcsrJEzgW2E8Bo07WRsxjWeQkjPbJTz47z
Fw93ax7Hr4vI6RjGVqGsTI/IjDKy6jpyQ8HEfYZX+jPUcVDjdnOLsvBtF8mI
n2QpisvGEwDQIIv4aq6zYJwgaecaXi05OyY8X1KT6TaOMIDh9VxA1Sa2iJah
BFNsqsxX/FrxGV0nDiRJO2e63uuQDdZPof3agGSV+cKy0N85JDegA9qSFSkl
f7BBqIGpaG8rxRxkd2xNT19xpvqJrJXbuzS3FaULTf/MtWORFkRHMCfvYCcI
zjGZbgojcab7vEzN4EekmC/QuEWD9jNKuWfwxwGhA6wzoGjKHzSDEUc6BHO1
+3CrwOXj26xBEZx4W8O25Kmz+B3KSJUl1lMykOp2FmMrfYA8AljkxOJWLiJu
kohRNwdZCt37S7EjkYnU3HScY6Ovmh5Smex8/sYl0zqySXoskvQDgLlq8Qh9
XKCEJL0TumVcUxd+yR/IrwaP9ZWQw8ymMU5e+kt/YHYobWSSU823630WYI4g
0Lm9R1UGTfhJrA29zyFeN1ZcA6cQfikQ74alFoPaEECFpxXpi4J0+PtdfyQB
BGUdaW2iZmfFnBvvlYKtYGIQkY7KaFRptEkrKDnwkcuYOfCKX7Dy7ceuJjU4
lZyRVqQRsZCsRMdkEetTEDzS1IgSSA16w1dCbtuLamWFfjToH4ncps+jb67j
lVyLNU2+HxkNVx4Ar/zWcWVX5wFOSCRHqJ6bDw/bIHdpwhoxVy3sMObeoXPf
otF8BCgMhRHaGBWRjyFwPJo9qQoZb5u978Za9VJ9i4POks5iq/LHXJgpuSSs
LTUnuyUx/eghe06KDLkU8tzL/xcDk1c0RxmkX3T+GG4VnWJ3S2of3oGwovg3
r0x56UXhaFXZSavy8H0XMb3Kvv1a0XSFPcX9/U2urdfykut15TikEIel3RIf
xs6EwnKa4uutX//QckYFtPfHLu1g6Pmw0gvj2ZGRkIwsIi8t4hWsFgJmZiSV
Mv6wbpjoNQNjMyZ82iK0o+6WFRHUJkAFGNQHEOoQHTBGqIkrI1BSoLqXSul4
G4suxUc+YrZcmlDsNwUKn9TCI6MNBZe+0tQQJFgnkEwfnvMpeK92f9I1NO6j
Tn/9ac+1hvX7IJiN0cNmpVZQ7BN0gx/ueCmkFEN7ktPM/ckrBg+dbQPEvT7u
kzUaa0x2j38Jk1dAY1kJpSCBgcKkLkP4mZIvSdkoW5aMCi7dYdI84zAOmeFE
HRv3PPeU1zhs08/jL8F7ipFBmBQwF18LR7gGnBtMB6K2clmUvw4UNhE8mfyS
Pm4JH7jxh00KNPYIYWSwGaIt1dxK9ddDjqRV/clDhvwfdCtGNrPfveJX9yMf
9bGS6FRiTPm57B3nAlUmiCIy7Iz1VdN6cRgevE9682W8zC+h+MamjSl96qgL
EnkiDsl5drs9a8KNH+I2ynxw1D4W0Hrju+ZdmYnQIrbBUAlFDRM7eYXtazjB
/Alg20DKFlBcbx7rkdp+iOsEjgiC1ABMqXAfqYUhva7+FMhOwTu1GiOnAxlS
QNOkINvwpy/xpDDr1DqYLrv7sc/8/5EJJvFQs/Dpwayr+K/aEPdKSu37rOzQ
yhQM7TtNTyXuMdaeSm/SUlZbeBpcmRFwFR5txviyjOXUllYYpRw6kFSndjib
90xNzluAbJkKkJTsLz7XVBdHIQWU2PI0B0R2yOWPl/BiELxwZQHLAQtAmO67
JU3kA27K2d1VZSNTYWMaexta+z8OiHOSM96rf/fZoOiBo2yY3DwjznN7okV8
CbLq2ByxkPzWicrdcQbNEO3sIojl80qPNxr7dw6uRy5KZRFSgsKvLwbBdyRP
cu2PlazFs2T/UPNgHbUvNCKu98yVrJ2kT7gEGEQMO9rd1X+PR9yz9/ukxxbh
XziqBN9MDdVljlpPmDpusV/Xwdrc/M+yXuJahn2mYZWsOjDZqVJWOPMIWKo2
pyBxF/Udrt3u32skw8kB2Yq1FSgiZMupqqaC68AFzIrsYY/gvlUzmYZtv326
RYAkuHd0Dm4CrROTvp3W/1NNranJ5/Ti5V9A+Txb2EaZ1fUijwhQtRiJVp7a
iD/7R1ytlxZFjZSSA1rwWbO5sg1gALWvcHFutH0RrB5/A8Gz2IISGfQ8kLRV
35DyK6ee7qIyOKQTUtzIvzIDs7MAmgWOf+KT3IzbhSXXxE2JnSCM8MOws3mn
LDl499XstULocbvG2ALvfCO7O2eAGl38CH54zufgeOPwquNCP+GnR5DSu/WM
PCO9MGUE47RaauZ9IBONF/HIXHRbplxqrerlp02yrKEdRxJQjVWOAN58qUaw
oU7h3sjNV1rnYBSVarSJDOyYYpri4s35hW4XhQR9AiMj6oEqrL2aedhdVVrQ
qEqLneGqg3NhuST7YP6ut3qEoMTi71YuTKFUDG9AU20HrykItK1zPcwNQLrF
nyOGuRpjap/MELT0YqB08UD8ZFBKJ1ifQ0n2+BenSyg5Cf7r/aqGyW+IzTE+
ElxtKbTKuJsUJ5IIe/bvOdhjcN0qUpI51vc/ggOhJ25OlHaBILV7NY0NUHPY
d5u2BvPNjKD1ElB+olfKedtEVKKg20VbY5yqbD4haGQZtt4KnP8vieUahOqc
SVJ2tQxVx44qdPJHduqaXt3Cn8R2nPChvQdOMIfG6OFm7Chu591cIie5UW5N
G22rqgG+mlX0tQkmS0LWKjnG3gdfC/gvyvP/EcCz8TwsYi2rSPRWvZId9P+q
zZNTA1IaU/qU3oQZM5htWyux0+dsJk5rZoGZL0bqnhD2PhZ/55XIiXmnPdNo
MVRf2Mro+khJI0qRTfqakuAOna5i6xs/lj1AGfH06gJV1ezrti58EH4ISSc4
WAoUr4LkLPjDcIjfKw2AdkeQI0BxmtEjTseKbKaRhwLHNw6wd4fj14PP73T0
sSvVjqTOjW3ZmwLlN0jPm5aCKrWvjgYE1zpeo/bjXKsYtL/gB/fy0tP/u3FV
oFqd4duQLy3fSi6HHsRKAUG+H5sHI6UggGdDRxlWDy2nTZhFoLT5FSdoZ7MI
smJZeo/K7bEQ6tDuJu0g71xEeTnFjMiMt7yppi9B+AejQeWedMkrCgg4JlvA
6lc5/Gp4UYWCtER8T90Xu6S2fpYBEQIdk4KTyrZ4HaHZauvo1gnqhI8u5APH
0DK4duGUjqJq2Ih8YQaemBTK0ElZ4Te2mv1ITuvR7Bw+rXuedJ2PuWPeQsCu
MOF62Jn4Vb5oWsyhw77duV9QnEIndwV2CQT9zi4w8YPqqBk3anNkb5D9Nimr
OMbSzIwe1HIhl1LYfRriQv/CeQyejjyQmh88xX6a+Clhr4HNabIOzc0dZ3y+
wbBHE8hCZrH/PncSo6RGBULd46yQ7ZF9K1jPmdQtP6WRF0VqjOa8rmw+H/+O
dRkm5jRv7QgZcnJVkiGKW0+F8XbL1BF/Du7bCF1IJ3hlqnNcb5fE3hNXAJB5
UYj7IFIcTpqmQ1JQ830pYePosqFKIPCeIqA3kiURdZwppILKGCsufSA5o0IX
GH7JaW3DvRcHNTk7YlY6eOG1TEWyNyU3e54qvIa8xEC0HqHG7Fp5eqG/BY40
dNeE+Jrnqkj7Zzt3srQGn3dQtKITjAOGqGKoK3HocFa/+p/+LoJjPU6mqlf9
22Ba1AsP86/5B77dT1DHYcK9rPup2GrvcB6s5HveqF3OgW7sWyaTyDNEumGq
bfcoFxfZLygQONUSiCz4o78BP16PE5TCey++naitoToJivipen1QpGcx009B
qpsmR8ca9pjrqJGwjPtM4xYJo8jmM4HY9iaj16yCob7KXyYpfRaUJJOVTxGL
GGeyatFMnrcV8PwHUc+6nbLXh6C8boITKdlK1aYgmjrzQzoujLdIlaSl6xT0
7mwYO9HPqJSfTbcJ5SBCt/iwwh5t9ZW+qRiso7XSkOQiX0wFrCkoXTy47lCD
dNcCe2F9+0HTXQvKbn4FR76xWlfLTAe5DPsAdbVOy9SvN5Trm/bW4MXYh/Or
Mc8EQqYG6Y7wsETWVfdxx9vmk65LAzuUXXOCMV5tKbHTIAhRAfppmkLMwROp
MgepCm8xjMh1Pdcu+1hfzXJWK1O0lAYY6QAJjPjAdSWNNjhAqCIGmJ4CzdJj
Rk2UAMUSpqchcSqItvueZtIFo3pYbfB0QSxkIc7sccvmfcTNH81GL38hhen4
dXAjWtTOQMImx8CGGxrMYeM0xcRT41Ia1+zvVYZseLEv8clgBFnob1KTMOBj
GT7VcslH7Pp+zMD4+vWYFVy+qITUPSMMLJHlBW0EAPWXbCMG7THVyY5+BEYn
ey4CSuwvOF8FTMNNznIi4zZWF39S3vcdGcI4G5jWzni/roEBaf2e0fYV9K37
QgFvd8jyiQO0lSXJa3jtnczkJWknskneB0fpC7MXIw2VhaitnBX0YZ0dlNBi
b++b+etoDpYNXSfX6JCIaCGD2AflVNGY5BMOMg7i6gC+A0/h20XI5gehZHZ+
WmnMEJkNDlRBnc6kSQ6TtvArkOfPCGsruYH4XIsOav93H3i1x/mh1gUmh3Kp
Q15NY7awHIElTjwCCUpgcU8vgd3iKJaSaEr9Sn5/8OKHc8n2Y4znGkM+1ipL
YNVgssh7etn7Mfc/KP5R5tQYOQGIwPeLKPiH97b9fun5bV65QTWeOWvdJKeO
zAIaFF1v5RUqfCihdlUe8IqA/3uHAENjE/D/npbJXpeMiqXGui70rnm5PAdS
QfGuTfNYvnci0waE9A0ULB4EpGCZ8YWDwpf9Xxq2GW361kLgmtHRPvfW8y74
SkkcR6ExkEJeHckNyg1CHP78uQn5e9Ly6wILplAAf51yu6Lb8rPQLx7LL/ea
LniO7DWDQdbeCoQo/SyBJaYVGsBTNLuNdzwgGylAXyq3JI4VNRMLSe1HeFsJ
mXLQsHUbAmS2EBAqwHNc26Jh75mo8wcuIakhWBv06mP/JJGEBTDxLMb/3aYc
cwUYVerlihy3Zg9v+fk78MIMgDWLzaEtQBjoXA5vyfO2Mt7v+p2oHWc0DLrv
d0n1dHsQdaGDeJuwNzx3E7a/tiG6ST3zDCb/AenETJPWAN7R2R0LAHLSeHNm
ZLe6VpvLm9DNgiE8K0IBnUy9X2L8P9/Jas1IQwZNkwe0IkvucGmetHz2VURr
W3zpdDeMw8L8F9pUej/1QTkocHJSNUTleV5pEmm+enQUbNy2yHT++bft65OO
b6d32UsgKzNNG6iwiSMZqInI/PzNlMen2hhY7dQSNG29P066gNX/M2caWaaF
t6KwC8t6aWBjbq2rr46XlzWFCe0PTbVTBGq8LcDIQdTgqg03mKHTVKmQHjlz
IRGQ8dV5bM/gr1buiBjcPD/BHC4/luUnPUbehhaMT8tm/aVF2MqA46hk1Oyc
ZiZKtR3p9vu2E4Rr5YgeW7wGkQL9U0A++fxrzWVMNkKU7OOHl5ZwVIrXE1OP
WKsAMbLEuLUK7Ox4Lh28BEjHq/5EX2SIChVY4Afq00bZO42AX3DYbDZQ0jDF
EtUFFOO9UQmSUyeRF1mwozOcQRKa5+bGzWfaDJpuVRSDtt0rNhRFcSrs27FH
OF5g0iZM/bHDIDUmuBPXnVS26fxT5H40NH805IjejlsIkvQwKp1Bdxva7fZH
0XcFay+VmDHHvz+JlQekAQa5oECJ50R1dOIzA5ARQ+C0ytfnZa1gNk29o/JQ
TCK/zMwxqFVNs586esruthsnDqVM790MnNE6aAeh29BcCoZOYa4iAe2Afirl
u5CgG74tPqYtRUFvb8HKfQ/SJVO1K/jfgQuXR/9K2s27bhguWhXH78+RyMob
iuV5J+r7Kwz6bPAxJwjpxPpMLCbmC3/1WI7DPvdYTiiRgMW87bgCxRH6oSkj
k9KitjQvpneLdgTnUceW3FEJS0wssxr5Hq9sB6JVXrtWJxl1ZLjVHCw39y13
rNtOWejGakiB4Ky+Wg/Wlcmh1Ms8I88Z5OecMghLm3jfoUPr5I7sUKhvRXRU
iTGWcx0KfRsp6WekkLeMmuBxIt3ctJsOnpBJ24CFWOPJkjCqaLI2iVfe3c2U
JI5HTvafuZQO4G3r7WUoFue76B6Q+s5z3+PXJE/WCZSZuULi1v6YV7lVj1QB
EhoiCzntZi8x2laowr/pjEdNnueDOYDVUTAA/vYqJBOH/FwvM9jw1o6iYaY9
qpAeVkWIEjYv5G7Hm7pLY7rmfgOeDgsDv3UtO1c/ISV4y0EyXmcjaWWIykTo
58Mpp17xsBK3uiEvcAqE8mqFM1Wc74fgdTEpDaqojkiNOMNrkKop6Nu+9/pY
gjiirYGLkhjjf2ysYt6763TKtgFmqegm9ne9Upouh4WpBsC5Bzo2jpcufhpa
vRQYESUHUtF7DVyaUvHySAnMq2bk1LZNgNacqI+59JhUylmkUM03pBpBMTOO
scPyuGIPUmqHU2RXterxiTcuKo+COiskhmZfor9kKr9+zsaf5cWZHpkE7Ql2
7c27im528cJrHtqFpi7rk/x1tq7XXb9lqpxjdWz7KxFWeqQOhF7s7zu912eC
sNsVn3Q7C3IChW0EOMQXICNbAL6iUZqBwzXveo7F4Y0omu+XZ0VheZQxQqcg
UJX9QSrEWy9+/iKb+szLqFbIbZJ/oURXVaIJbAzpQU+IpVh6kaHVNj5LS6Qa
x2EaF+f7zNT5bIOvla8gQ3bIYSZ5QFX9kumJzLEm2k5Y8LGOK06gdF56A8+n
e8TOi5WTUWn9DXihgHhhxwh7PhTvVz3on5rk47XL1ZJDov5mPWpV2z+XZG4x
FOJ5PZbs47SQlWX4Fk0CJW5nhZXiRhtDNgdvl9e9Pvg3Mwit6CqYH6tXm2Yl
lIE/laoUyvQ4qVmtlFp7vHcvnKrS71LOKP1YcI33WY76Ue4N9HUqQL2xXqg2
5jOjjAPF6RNszMRChl1P58O2mzvPZmJTi7pMThm9a7P84vKCgf2/pemZXqjy
dmI96Y60Jcqa8iXn90mZ/YTBvdvbWALoPDdYY5dMCRROcU4kZ1e0tGawLKQd
9Yu6rhBNG/bm94LwqWChb0hFYHAs/GSMs3Ez2sdTYySxux0FngSpCHXysxuE
FrcWV3TDOwluKGg8eQDVCA3uxizL724130anXLSIePI90G7aJxzlnHx4JydD
mRZUpq1tjDvQIbdHPSTXp0Ci1CYIxcamRcEolZHonktsyUUaB6bQQ/D3e2xG
+75QbFqfjekDs6lyuGcApX/iHYxCAwP+9NrxW1q2G61rCS/uTilUXfdHYSuG
ukTJnxm9n5W+f5Hbr4DT51ky5YBDVDpxaPeIpt2ZNB6sklIxytOuhN5tn2OJ
NBUIjhZbSHtLQD7WiHTas5EX72MLQbtVqKVgR+qNpipeq3LaRwDDGePnLq9y
zOd13F4rPGlQYxcVNmnxrmWgVYDCw+UO9DuOC2m8XsSzV4SKSeRrQ8NdIswJ
GnfVwOvAuYT/SxdwWSqi3SdYArvM6cN6lSFAPigLrvv1GKfuufBPg5ZF8yY+
G1EFy1s6qM6d/SB4GbaBY33CIgAd2txQsq3DASWmxXqNnGblx5ZVgqkNPenT
3qAU609lGseDl/7FqrmIplXXzBRG2INemxQ5s8VkBfQsx3vPoxHRUQ0DInJv
9tHJmzBdCGJsibWXUnvSbqDtESDQ9TXgfahY2dc94jT/1sa4MzZd+nKOQ0EK
zeoF+rZJ3yROXmVZcuVwTnuDkVGZLVWAU+D/GhsCPOGs9QQPqZnGtlofLyHh
DnNZOqMIVblzIG3QDVARXEfGymTzfDkf8/VnKNBRSi0cSwCd96q/rzLhhEbQ
dueW1eFrgGfOOGLcbG+tJVHFgvkVXCPWwHWOGUdXOHyv5qmX9t5KeTZQ6+Qg
o3dtUTege1ac5W5czxlesooAuxkL4cSpjaMBBN/MVQBHohn5zWY+vi0vqrMg
MOqDgUoSuDNkmnLc9M7LKNDec7ukoEh82dVV5L7KW2db5dKN5cjvJ8UHKaJK
5/BzsIZpx69gfS4M4v6JM6SWDiBgwb5+rZVgodRYipltmgb8cZx1e7AXs4cy
fylLEWtR5OTO/M1nQ68ZVW6LctdxlSlrd7qs0Kwmp3r8n4446SdlxE74Vc5f
r4bIkInMGtKZw1AXNQM9ZWxB2bBq1e9PAY+LQOn8TZWsAhFtpP1Ou0/cmrbh
dI2jX8a55CyqkoOpizgiLlJV2j+UVxtA4WTTFufNiCD4UKFljJ0HOIrVOEGM
CIfw8OtWkHBHpUxV9oktSIqMzWMWHkuE9Iy8oguucgTUp+9nNcDYRUkfj1Zl
ZXhSgbUrONp0VPqOB/90QnlUY2eLjx/9R1NfALFs98dl3R2FyYyEHtopFJLM
uNQ2q+Ld8YfwFgb4HXGIB3XrLagNyeoxI69/N5gwryIwfXp6EvlK0uXw+Wts
HtSNowt1gvlKT9CaD75g3hh7B6UHkNTgvVmmsagIbRKB/NB8eoMrEKweSs9J
FYGPtMK9rrgdnCKXNYKLgAmnXUYC1q9tKJ473CcSbel+xWqlquW1+3cmL5Ls
hjLTdAVjA8Ib9VgMHf2ATDN1r/obVxfHf4VpOR/REQFTzJQDbuErPoo5TCRh
WzjEVq9WQ3CUYwIUQM/pSQBxjzSLHr8mSQKWd2rvxocsM655xnZQ9zgRIeYJ
iNW/pvNK4432IsVfCJNMJYhLE3Ejb1DQZGSO/Z2Ie1qj3+cbo7Zb2Ny4ByUa
IYGvx1D9oSxHfPsLX3ZwI/RXM5RKOrU2itDuJ3GxFegZT//vwWGDiUoFN7gf
lsRtsjHyAtVks1p6md/CD2uBCnX6SPlk8yFwg+YyT1lTQMf4Dy1jvCx52iPF
VmWDvl0Jce6dgeRdttw9PrGWoSCcYm7F3yNRUlD0RlN6Zql8Ta7Lazgx89bi
Dnj7r6ePuOK1Yyr4wi6K5GkRz0yAAr+cUhQR9l59eo5C3BZdvc1iCZ92HTGR
P65VBNvn8A/99XS+B/5dAo+BvPGzBGsEhGP7s2yzBhkLIUxhGEvlVYWGIMOS
SmZwk+lPeoHSlQmHsskmCugU1B/Z8Y6LulAEjNuhII+qRNCXU5itZ1+9qfYE
W4auVaQGWIp5swEWJBllsb+D9nrvLy8LYKhv0eJxGD4uGItuo1doWP+KmBmW
oMau8/9RMkoOGiDEbhoeY8f8Vex8E77j1ONcKpiSAtBec0swTueMDyatd/7o
GN95yXNUdO66vgIrUpg/qSDVVygGtsftnY/WrX1C/dlwDf4NwqgDXOD+rjp+
VcfWYSLR82edV8e3ad7/F7CSjAlTarsUuLUrw5FJo7ItkT6IzcD+OckG6OKy
WffsnephehYpDHNoylPrCsgC1h1OAv40WiE53RkW/UZARWZ/FDcOQWIqlrin
5fJdwont4wR5fTKgQV2tdHgkRSmEosPpBCoEmWRW+WOvy8FxrqmEVVMlWEGk
Xsom83lfhxHskPIwCtGAwcv6U5cKmYQyRj8CTKTgFGPXYvW+tPtIVqLY7uWe
ZjkDQB/GOoynD9Enw+2smcrXbNCQ6pBj/8C3UhUZ1Dk1beJJu5Y+I/0uJa9f
ci4Hf+zTZJNADExo3175T4W1SCrx7T2b0MfBEjj19e3stm7+tBuYUUOIluXs
GOzz9ps8KkuMbKfcylUbU1ugmK5G3GKvxv+LKCyyJ6571rshe+dsl2R3wkum
mrNi3pPatSoVHTO3POsxQWeo9uqWZRZ6f+R4jhKrXT9ATUdQ750q2DAZxtuD
1AT1Iaztpqo54T+tnqrcvL1+NL01Czap8pHAYlie+7tiwtxyZfpDxXasB5nF
f0vuJc3d8wlnZK6DCqKvrPryAe9Ne2vuZvKHyQsQft+0gH4iq0rx5evKtFzf
hXLdBJKIgSKA6lWkzmWFqs2hzjkwZuYiTVyZ8eKSu5qSV7qjkyWvdSKYS0Rk
hl2CvBpNcMQ/BwD1D7V22Wf9Bf+6prUYx2w8axSVQxVkt5PZ3qHkS+4mZI05
Hk40u71yU0rV5cBcuo/T9+6bN5l8T7NfYCuMnM1r48CwyQAwRl8WJ6Vg0Jn/
6ivr3plui5lSRbr7u/b7WLmsk052lCLrHN3RDNF2QLeglSJ+rLY0jtQGQimj
HpuZaHJn9qOPKBmgMEcXjCA4FgRVoBFqaZ70XAaf0JwS5s+cwCSRCw/+ZZEW
3eEUu0kn+SpWcKi3JYiSM+JE/GQ/Jhs1HvZL9XmCBZ74eQU01Qa7K2DkyiZI
u2QgpIilJy9t5uimJprMZ4MLjxEuzkt12Nj7wwn+7mH/hmejry+1R+NB2ESk
1eQAk9D1anDZXwSxAQZNMyKVnoPgRnejT2GJjjpeZl8qbjMg7y68Hn6ocHvV
OGm3h4JTWdl2zd7Ra+cdmkkFPm/V4drRWCJKnuRtlgzLyscxcvNcJRyPfMFD
o1ykrrtrqTT4MD9rr0msoWF3l1q849De78j6XppW0Aszq3Ic8R+3gy33qoV8
j2IChZXu2cOQQgxhOlchK8J0Z8R+BzGxNViCj6hlPUzROaPCa9TCw7i0LpZh
K0X5sXkBDcJ1Y78/Vau6+ojM3gLqbZmr5Uu7A9nyF/uONdz9OXlZ92bSuYMg
KuM7xZxRnK4gUFroEavdqhvyijbLoDzzRKSHmThe17uMP4xI1KRAb8K48yer
mg/WFTo8dMVf7xshWf0ZhJeJANnfE8VMxK9LV68cFr6fMnGgcYKsdoM9ZmkC
w5SierFOEKfN0Yp8Mer/23BPPrH3lSvV77WzGP+ukWW25HxbRh0PPekadD+V
fo7jQA6zIDbvNKRpI1LjGr8FHQ20FBNxLljbsV27gMcyAVqBD4cqpFfyzqPc
K2o/tEgkCgpEzjHw0CsePLmKet0630k+/afjPAcS/FejPhLZTZ7Ea/28HGfs
Encm6pMhSySiwndKfXECl847oGmbZLqZfOkxn6Li+mwaT82fPVcDmD2kFyWc
z8j/6mbWq2P2Bj8JIT8UHnwd2CDzEVNq1If+bbsB0XFSkOlq+pdqnRdLS0Y3
H6RoKUvoLz942rHwqaJhmc9GEXcmqfYzvGmi9+1R+MzaL/WQQo5+kscjCKOJ
oxw0/MsE07B+XG12bpUNsaUY/sZSYFo3WjAxvoH/gnteyS663/ukJndvcDqN
wjI1OTI0XTY0Oz5ajQp5VOtcA0y8GUOTtdrbjjbnQMsRLKkx0L+4Qil2TrM5
2ackWrGobZvZdHmHIBMao0K1T+C81iJ81RhvyFP6er+4tBXod2hXPMnWZJt8
puoWPDHaMKu0pdDKnezlgOxULxgfK8pDvbw041StCnm0sKkwIJ3CGMbwiBBg
nr9XRywULQwmUJfTti4BbVVVGS7daYKSsEaokZ0/XmXs8qTnNEg209fOHv6E
iEcMojt/WACY706Mbkk9mv+ONmAHxfjojOLXtDIcTp/iNWAIAZybLvuGgjgd
/7Fkt4QdhLGO3oYcxYCkzkFIBQoeDVNdWCSGuCzGfu0YOYMPAdmKd+NlZZqg
X+nmlEJP0zMFhqNkAhf7/+cQN8QzvfU+l1qd8NGXpggKyMdHLNqVIn+3e6Qg
Ggci05H/eR74tzfa7DsydgB04YS50JH9Mx+lJz/TsEI3P4+Jpfzwdy4mcy+6
vHBAv+AdYYtBTAx3k9qCoYZktYoMPzdNf9JXMwER0HUUMcOLNUXA8EdgR52v
JLFl6Z6/Eo4htLy0B6yiYNcsemZe6aHimuV8Eqd0YneTHHs1r4WXye20XhFB
uzzQT3Gahrh2j4eu5wIWZmUZrW46ofwiUjxlBu68z5xVDaMi2h2CkrWwDxqq
OyyQTmxppeVBQw/FEnvtGx+7b0fIg4RTu8PgYu2uc1vOISQ2rXNMHYki+93I
B5F+ApCcYcDBsHdXxBS9c0kV3rj3NTmJKNkoRKsFb5o3Z38swtZOXEPNB2Oe
rXX+Nd/BQl1yoaiifCfTcdPhJz/APazwpQAqDyZQZlaLhObJ5Ro/VZkXjMZo
8Tz6zGdnjMPuQ2ABGXif9cWYy4t3ZiQyPCMcD0sXg9Jw6F3qQG20+dHkdWxz
6Kfr1HDK+42l54eT+a5sloXQZmGD0/ygZ4TtgZdK3iUKteFQt6WOUhhn9bFr
HEwjUsp3c0WVP5nNfCc7O4+Qcq+w5nQ9CcR0VuWMy+wpTT8JwntnyseqSnnO
kr1gPL37kohlh/xMxC8RSpBOcT7A1Hs0Wx9DrpwBQtFX1zdC3uzNtZ3/7nJR
hGqmxNNgiok7mPc2lkshelQoFl8VgssyoHUhvMHt4sB8UUTMduMKrF8QXpzZ
blhNofHWpzewgAPCu8RGqXgIQfb3sZHMYcuO8DfA4ABkZz/0ivdfzvCI5dVP
55I11GwVfvRcMIPBULhCzKrVew5PhIaL81gnIHE+PnoH696xbfD2Be6jFhuR
BNLU8ynSodg8C3sZ/x8/kN8niDIngy0kiGxSaqftgUjp0wAeg/vTcjnQKE+r
YHKgpI9Rh1ycDin/4WAtY1rNzIbXN82CDLAedB/AwVnpo5ZpBBYiJj/6jS+p
VAqDNLJu5gXw/73o1Os59Uhl77qKu+zj1WZccVf/BKXFdE4Q63UkYihuvV6y
U5qu4nDhLp4zxiQ76DjQoDU4yCZpHdl+hj/y7Zj2HmVKK3uxRg3Sr6hC+kUn
86uCCpQPbOHbTW6Pc2FPimcyRaY3ij367h/H1BPXl5fTdOXISvEr0tZ136sH
BasIf695LvaBaSKEWzUiYKSOc9c1XLPlLF/maCudCqwVS8QQJ3pO1TZQOKKG
fgEMs3XQj7L3C3SNS+jU1bzQUwQg+IYWrZTiPKOpH4ikA/n3KfkLtHuF/kxB
dqTy+YU+MXfDYaDSuFbw89JsQcn9RfhBal+SVXb2Pt1HsMIU4zzwUnKLMn+Q
QUxerNPSzIuG05XDsTj8Qg5UnpRrLoLMvdrOJJqMXoafvA5T9BJJk+Rfu/o3
JlRtXxP/IPKsB69w4KGdas8fE4I4KVB6U4lk2kllK5RWqKPf57tI6oIjPg39
swcOcNQRQdd9ED6sMx1H2WKq/GgXEXZBTIpEpwCUBqUNVEFhVVOeS6VBE1CW
Q34T15nIfp5F3dwsgs4tF1+QcIw1y92ChBoYbciN8xPTWlX3HmTAPIfm6j4t
iZIh5d7o/ZQcrPzPOFRNmcMQHosO/6CRQWuwqv3AwdwMzZW8yncAjTgK65q0
W+dQplKYUFGpJzjCXpB8M48yb2nVPR9CqRav/I2zN5SVVyFvkYT/DIlTLiIb
6yYolMbkNaB98Xg/m1WcQIagwutOgc/tLrt+Kp2Qn59sQDilY4MmKx7weVn6
6aufh5jZ2NGMQ182c/zHczpeMQ9upsXMZ+ciCir2z62oljZVIhmn+Nz9b1Gg
NavjOM+0zeVqvUw4UTIn/MTIY2kAtesMlky5610++gm3IlM/W2Rc4PomQvx8
vk5CfgrARRDRCI/6Wrp6lG7f/i72wpzMAv+JBoG/IJkJb2jDCTdGX0f8xLcL
T7tIIH4o/Oyh9u0F7+35y8quRYdkXHxMUOf8RynKRQxBtUj5eZe/h/PM30MS
8l2qi7e6Kg/E0Zuo4Z9f5QfbJDUwxMvsTbI7DgnJj/dADzBSBRquh1vWxtFV
tbjkIvXhAZ1t0/TlXFt8cRFR9+LidKOfpVcpwE4Ws0sG4KIFjxaIHPSX/5zJ
Xtbr7bXFNukUgEilpi3HeH5m2LKWmmEVlhoyl9KGeNROj/SQ/9HITQgSpzE1
o13CQHT0071v9KepcO0UPoWkkh8Ak8MT+9mgOMdN5LTr8FIkbnLxpogMrfyb
a9GyO/mykneL359LBAQ+QrmpnC4FjAiveWZDkPVk4ECwiUYIH9jsyi9XRHZl
a4oxj3GXvPXqAiZR/hKR571mPqs+qvCBDtO3Xu6xyBryMvJQ4VBx60CB9fOK
NZ7feVa1gcDJUqJFcHHBlp9MxMMGYSRukFsvg3NCI2D2evJbn/4KmUm3wpDi
o6XZ6jnRibP1OsPIjAgFBJ/RHJxAVeJ1jyTN4otDM38LtGuDgTXBzH9R2rgi
7U6wfmnnWkx9KX3Cf4IW6jo1lkLaT+YXV8veV59gc/yNkOrl39Igj/U24ijx
D7cJw/q2Jht6govIh31wnC0jYoQVCMVGIntHhTMjF7rh7q23CFuLrnbl2EKb
/U9uGqeQUcWgiDKgB5BYzlsqV8PV0EnPeuoSLzcGP00fdxeZC8AgwM2pjx7z
C+a6nZBhypJC4rrL6L2wMyTKnBEe7ovxyhKp1gaIDB7Vn1StML2bHUxHJzlw
EEtxlVWsHM8gAwenXTeNYMEN3fg+QHxT1Op7jz7EwuiV13ZRt935tMl9xSXS
A/HAxmiX8iPvfdTr7y05i58vMG0arzBnYv3ZlZbCLcxPvLKixJm9IiE+NP7N
vTZ0yh06mrHzVIaEkh9bd5Dd/0ufawSe5JHHRHoAtuPUT7wzkQ7aAetRCYDK
JNn4RpBNA91N6uqInMWB0MYMPCYWY9+YsppWpbdrlp22Xe2ugKGr8VGsLoaU
cU+OEXRJ4VvqZVLbv+Xl6V6z/T1MjYR4wUxMy0II+xADMq1qBx810YKPL9uz
UnF5z4WMm2eKvOFEeV3hTXs7MW7WEhHtq7H2YcuiSuuEcZm9BUkRg3CKGu7Y
FxvB86mzcMaEchbLDjSs6CNjfpXPw6gEaotxFVW1mHBJpFofdFXn8SUO0331
9DLjA5nX+7nAfUzBHRy5UCpFvslWsf/dbIyrrdFsStc3or2iz2VXHs7GGvhl
1wx3YrdJpuLWSJG/+07jlknQeWof9KwHJZHWtMw+Nc3+Znzk4AZ04kwee+l0
wizql7Kue97uJmCOoL63gS10LBgS9Hw8EtBFxOAIAtRiX3R8+epPoQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "5PBMlWQgil6yX8ouZKsBn4gxG9o9nvffJEfq9nnkQpGeF73RhKsVD7WpI6IruH66K2SowMQUm+mhxDum1nApCopr7UehE6NYtkPlsjvVBO8EWNdp5H/tcSMYD9anK92MEWl+XfvD9rPEAuy8rJDU2H9nywBUht4ZwOjJ7Gdk4X0g8FfTi1+/kYeZrVU9PO1v30/4O2cImn83Fkn1gCW9sFNphOgexpeRo7j9twx46y4Iarb73b3+5HddT0ZVbZVkuHbOaGcYaNlk8TAN8Ix+Tea8hSgjNoet9nyF6976jLO1ErVcCxZf9CGcQPraUdApNMPA3EiKGf6zkfmI7dWTXy1EhVnEK1bV5wiu3m+zEp33ObwYOpHxynT22Ja1X3nb3oV+b2wKa2LfEi4Oxd+F19EK087qPYNK8HkrHMEnLOvjMZtfwjn1JyLzaOPjQ/WiGh5TaDPDx0fgQekb4rc/1Eg5e3tE+DX8wOMxvzxQn/PWKRA3oPZ7vLWSD3PVzy+2OfMWmrabFsCPiobyBP0Ut2vM+f7FtjCZu2lErryt7/fQER1RO8Bkb+YhWrW3tRLchpOgw46UniFbrbiWMWn4hXTSdFNJm3uUdSUOeZn9lRdhvWa5uOioNo0v/EUPCxuT5PmrTZ7wY/51t/b8g4pLpE6j4w9J7IMgjeE+u0wT/33NaC9vPeDkjuryHV+qec+OoEHTMyhsnSR4snV4SUR6JU8Yo6gBnQvKjOfJKjh+TdC7BAFUgs2Se3FgMhF3WSs5MezpDabNkHckXQzUwSuWMr/mr7lEkzYU0A9bScpmb17vMdOsxS+pMB1/Tyx6ohtEEvVqm2apKqLro+cBLHzGS/gWUYde8jvRZZbynFlFDtYzvPvtbFzhlCB2AA8n4Y7nRIaxKlY5IRYfEa/pCdh8axo8EJSjCFO2fCG35ycgL633qmZf6tCya9dMhgtcc3wL4LEyFbreL4aeJ0LDUxWGkOpKQLe1ITrYvkjH19uR/0z/QEsf/WWQ8P9vD80rvo7I"
`endif
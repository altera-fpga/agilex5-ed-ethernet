//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rmSHfyuyqT7Oj1wo2Bx4MWg5cs0fQOMRFDl+mdfJE9wGI7L4+4I+mLkGRM0D
xSqal8IU3GG85cgmIe205AZSqqG/QadP8lrQfReu9uMz9caFH0z2t4RSDcup
jgDos1LJAZ5K3BnRoyBVNGXJEoiWx75Etzo/9lYxEPecqjJhkTsZ5O++9it0
HgCqNeRil2ZnxtBdtQ9XjQE/P14FeGBwsG/dXCHcej7Dm9hoHfRLjjRwl0qi
nMve80QqbIZJlqM72OTX7mVms4snfUg/JLet616aAm3u1y++5THba/DM6NaS
RrDm1W/gfCWqpZzZCbfd7kpMrEa47NhF+27Hd7ZYHA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KBLgQRIwDppOEZfsqBVL6kkotWBZCD/tYullhcLj5bDZACgXNYmymYMEsS9Y
xg4iZCgIp8QXburEV5UAAeqJJxczU0sp8AWczZxTA0Rl6lRlbsLD7Kxa4Nlc
I3De9Zg4M5ghqXSh7KF0hkJGaLiP59drJovfP84BOsI7C7qgG5AQWh3oG0Fb
HmBRLQ1CZ/DGrJoly7x7Lx8LWdaQShpDDyjP9dJEgCphf3X1OdXyY1ZPvzQS
GKNWL+8uQNbOJDQ42qIL095cGO330ZkeRchbjpzIjXV+FGKA4LuGs43nvjVU
eyl+cNOGCdioeAJSHVNSMaENLC08HmYIn54NiDWABQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kbE/UN191V3DLhSnbpxYVWRL+Cv/Xzdv4A5I9zwPcxaclXcHEB8Ku0EzMqoD
U6KMxNHrOx3GqpSuZ/z3YXrZJ0yX/rJBj+hg4Au/ddqUyVVKH6P5ZcRTiAXS
4NPMYFB0CXxyJ1NucbdFb8c4GKZhfUAUyIhY0zGN6q3G32WjPtTkvq4BE2wP
IuUaX4W4YCeeCuJGcofzyJGL52uyDNCQhrfLJsiRNfkR2FVeJCzYPhZRemaA
w2bPZwERPKGmDXcZZYT2mB0WbqxZyG5IH4kyqvuRmDCQtsqkypXQVjaOUo8Z
S/mxnbl3ovA6Vo+gnDdjYPuDLowtPoTYzicfV98r6Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hxiMNeOXLCQnm208ycNKteJImKYEKRUDuHvz6XH1E/swAKWV9ePyv3Ox20k1
rCDAj+/mNG0OVKFFWW7IlhGc9JpGGdFaMds81QyKJAP6SWvvcuYE7yA2Wevm
LbN5KYgGa14LA6vQZCZ6UZ8oisIHBA0YFikW5/xGWkm5dyL1F2UqBCIKSAK9
f58/Oq54q2Ct7wSWsztJyaHZkb01yZG6ke8ipUWLXBvxrwatHIYp+g4eqKgq
5siZI5hpJexFLypiumJZRH60Ykxtm03iYtDdstcs4Qvq6QU/LVLBxisTuygv
Se3zAla/8+vKbOo8SyCA/a3gwc63At1/Xx/qoxyUYw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hTG28BY/FrjscJtcALhgnLc1kEZIGAMd+had2tRelZLrYkHvOcqavWgQ60YR
AJiLOof8EWJgkL0PQ//aMC3RYMaaIXVQnQUS5VAY59AWEfMi64lYccLy11XH
K8KjtKMOOHdHXAevOi77ahSGuLBfSXztCJPLtWDjBO0ni4wa+NY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
P1uMcX3/slZ0EkPnWAnxlAGBhDyvI8e0WrVc+nOx74AuPJoPPweHrKCeUkt6
TlsuWEqU+lBAcpP2xeH3tt4a6ETEfE6UJu4wzi5fUQIVdQjfTpQXqezm1zlg
bNii71/qXyY9qZ3b0uxfktIHWg+IbRD/y29LKeYLuhQ6yA7/Cg8pvWwCBTZ+
I4NAZ5cFug6cZaOCwYmu7/QNDWuyN2QF1G+ssIWu14EB8suNbZarnbnhRrj0
mc/tvu9ZP8vuYLorfrVR37eu9AS3y5hbq4gY7UyNJbIKxIVlds40ezjBq9A3
4MtQpbFT17h20AlF8bu3w8ay/x8zbBmMSDKZXfctlyvbQoRoNZjx304cGIvY
6iH9sSrJuWrL1WHbX5blY63REXDhX6op/pFW3BGWE+F3H+XWZKVzWCQdDioS
NgM1EjGoC6C5siAjzMjnTTyE/reoslhS/dXF8tTOdMbFzITyLMtKAmXS8SbZ
ItxOiomEsvple++DydMEpxUsXgGhzfdQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qMEIMShtpfunWih6zLC/FmGbdB9whDxYFAcZe3bgiAmvtoEOnAS4snZw+qFY
ahIa12XOrNqBQ+CKG4dQciRwYbJRJ8GW0GPrLd7vcn2M8/QlxNcF5crDTAHZ
lotkWH12TcQ6zdN/BRzsUPcmBjLVcLWUbpNFqH1tf8QkZ297YpM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dEXcbBggAwMpJknaC8B7f/cF9Vx387gmVbvp3ZgLjS/Mhtcejvkxea1WW3tZ
y91GxnqwTkzPJqD9PU3phi0pMZFSn+asPjQZ7G5CRF1bD2+Xb20IKgSPsc/u
O8F6dS5YCLK+SKHVPOcZWQ/1Ywreyvb3lLm3Hy7BTN+tGEOsSqc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
l8IvTI3Cb8Z+oAdEHouU7icjpEe8KhH9G+89Y7lJYPrraqTVUsmN77zdIOHj
T0SObJ6oAEhNzkqZRP7ene5U+iAEfUABYwtMbuvz/GkpJjmjD9ZUzJoRFSn6
pY17vJg9rr/Mb789ayFqcL6RN8ZBsk8GAJq9OAECSASkGXnUTfCD87jBqCzK
BlhVObGk3eRMMqepz43V/leI382lRs7nCQErpD3kTxw9TTlDcrn8rGdKqVzc
JoSFBHprRTlhWSN96zDAIaQ2pyhTILrtWTER6Mk0555b04J8WvmI5YjfQjee
dvACZNuZPJLOWutnQYGK1+tHfxsz4rV8BRJBjCRCqyafXj2PVMvEqSHW512Y
IcDaDTTjjGWyiyNpmU41705Ny/QmBbmWYDtPS2vQAbhrRvlOu4N7oDTdR2mH
jc2N7/nKrJXHYRY6XryQI9htFPPC+WIZDEizFemgdZFZpAlyYBM5JMYV3gxL
zq/YWorA2bpVhKNsLYGZYO033XbY201h4oO96sf78tXHm2Ae9R1JBRTNJmpE
bhCfdaehOoVZqkGIuZ/ywVIxFD0O3+gy3Q/St0ds0DVcXlHQCCrZkp57HMeT
eysDLIecb9EG5FnnQhX7d9OXQpyop9GMI8aDOA7mhTXzjQhiRAXO8VJ2PN1R
RTUtxXXXtkN2VHCDgws3KMtPHq0AouvPYLDRzz5c4JItat8OOJmqesvw/ov1
Ha8YWbaIv7Kzj4To4isKtE29mhZhVPMcwHvLaB4KHR0h6Ccbs/DTGz1RC/Uc
89r+XH+3Erqg3OPUgqfCEoHGO585oYXCFt1Ww4Bu4Z3wJ4nx9X5cyQ5EOrs3
Emmz7/VnwtY824nF5skMdQQdr4gHToT5NUsGh1k/S+n0YHpxoccRIjwCBKL5
HpivvePCGoOXeBRUNr9IuQ89/Bq5UrQOgQz78jqNIYeb2meRG+0JK4X104pJ
0LHAYvp2RG32RIE6d7qVSIAaSaJsQGYLF/VSXh/K4Dv4oo3J/2vck0zHfwx0
TmMfz7hRzB54Dl7hNQNDmXqQWm5458lgBZRGbDJe1Z+YPAxiSr7xBPXygBZe
TzK9gJDOPdyQSqhqbc2QiHYvBYm4jCw473Xzm7L1uYes5gdaIhs9nGjqjFZg
LDiL5W0Jx4ysD5TSZq4HDrla7nGZIQDPACo2NhUPBwmvdHQDb0H/bvam54Fn
V54m2n0bdx2nL7+qqqJReFGymHxbXMk+s6rsHg/CL3Vtrem0XrpEJdccQgY5
5qT8QwO/qcxdoCbq4XGy2kig0HbQ+xnwqAotp4c7PqVdvKdOeqasD9yYlqyX
Cul2HXc1pXjpooTrr7sELk+VBPRn9pH3tStEUb+/f24A2t4EyHYM1m5W+rcD
IA6+XQ3k8eO1u9kJMAzMlYC+nxn7k5wKOxDfRMKfkCseDeKTG1qrg/c5DbUr
eSlviNJUmcWKQxZ9FnTADiX+Og87Bi7hPMWSG0SlTn/JhE0gT1ST1NazaGve
roVvx/vFJNtddX8J78mJBkzFuG6xtMTtl0hKWYwNEu5okJK+pRlEu31RCoDV
37sHorZJH/SFcBEt8djjONiaNs58x7815Huetq0JheN+LYMn9iefj/2WVTjh
lYiSMGocNx2739ohpiSAGo1B17aUsyKwlXlKvR5gsGA9OSGJbWLOpcw5R23c
ksvBcxiVHrq7ILW5wNissQVqGNw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI1r/nPknGPrCzUANTwEw6tutPcrfZGK4aK1EC7JAFY39ze2YJ6fAJJnQ/K3LQAw4+S9yZsDZsoza/pVq+3Y/WvGO1sqNaBuZ97pCJRmJTr+d7AXhgcForFuH51/eDKL3ZN6ISiMo4abjhF5TTvZmwhu4n5BPjEo6a/NQ4KJed4yeAKNEDEhs1Ax4CSlOvsJe/d1EllEMwdkTm2Ss6Nt1+q2B1VaP0nMtLzGwI4lkrCgPrHqiZvLAClY/ls7mzBzuZK9+2DgDtB94fBVR8AAH2Z6TzV7Nthbo3lYNsSIiI7wSOuvQqnZRU/D50mofTwmtV1eGcxy2cM56q0gpd/qJWXvkEYFiwpm13zJ36uZyQnZ8lOPt6pNfd6tzjnk1bspsVWoi93nyvtp/sn25De2nW6dLJxYqVmgaA3LcrM70wsrL788das7xBY/s6XgIJbtWWN4J3NuCdxWeGqkywW0XhF1KjFtjmueE+GoxnVF4epZeG11oFDIKuOGqS6wPBW5fEdX9mK2xjYjaLoUxla8/y9i1LtERDLUmURi1qsUCysq37oGVsi9K6FQBpU1i7lOfCvdDpWdaIawciapBifDkwRT0SId2lqg0gFM+WqOz30dJcjCdYUWNx2EhY3aR4d/HebWUIXs7WQ7jCYi9R3g7AYIkpxH3nFJWWBl8wuGqRrTjoOo/qysOx/2Z7auj6x2LDdTTobxujN0lnHShwPRmTD5EISizNjL7RPdG15jsMSf7QPSphDoSq/QhoIb5bx+Efx1XPJo2QKWhYYlpCey1Pih"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jEZmeh07qpsoTA+8ox9+tkc4tQQrqfo8Ct8UZAdlR0+kia5Q8eTW5HRflP/K
bKg393L6M0WtIklk+z8MJKpHAHYxFOHUi0EXQ5j3jDMXpzNeaeJHtkAS8WBd
fJbevV9vbw6/8corNLh74Iir3CnwK/Wl0to5oQkfZ/3b05F1Un0pIuulyUy4
9KVXvXoQN6GGZucMtRC4E6BLcuQmZtJiHhPagk3N9DtmjGF4B+wcYrP5DGk0
Iu0p99mNOwZ20OUlg9nbMnqXXo206hxgp7yk6EQHvZbjSfyZ9Eg4ON66WqzO
Qqbb+qXN00tP6+5kxIpRbBD9oPrt7KM5s00fF2xBhg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
glPflxI2rgbuyPmj1ouQ2YlLS2zVl0apoo1nYirgJMDIa8Du9/BWS/ht/N47
nV5GUlF7/lT2lkAl3azQHCyaz5t/OxX7Tyfbf7keB1OogFQPJP6ft0KgjzmW
fegfpUtFut5ON144VBQToi08bjlqp8lUP7jw1oMhqg/PHuKW0pZ5eXOC+ai1
OLPvbKUlJYRVqDdO4K81IBdK05M3zRriRzyjOFC4u72K6ONqRAYdSecJB67F
1Ayo6xpfgXrjjXlHyTOq2yg9gSkT1jrVWZtIpnIRPEcRWZVsVWTy8cKZhWxD
gzYxuAm674nseydxXw8jCgiENyJpXOm6ARDvnTt6FA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tCa5uGybnnlI2YmsFTvDjEygQycR2VIh5BtIeCsB2IW45SO6eRuXRIZTZuhU
p91N69xolZJqUyGmALbzS+9iQasJKZ7beAV/G/Wi5aR29N+85YzdGI4z7aU7
BD0BlT/qKotHDBq+Ke1f+JzOwc7WtJmN9E48eHzasKHKhaPIULps74S1ZUw0
+I0u7rXfOFxFELHEMGRJhPXFloesjPJaJjLuNx0VarGWEigvaxRDidTgXiuU
R3RF4vJYBxO1LOcCNM5BJ+K7cbwAFkKwy/w1QmgGPHG27A3g1ILZjMtQbrJ+
BiEdxukH2sbTd0hqPHqJBdJuMQhDvxpl9mWhbLTlbQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XIA1zHwUOWiO56XhANjISoE3rD3qKWzWcnuKe7StH/CTcXgdXwJ2tKW6rFzd
T0tw0Hw5sQ/NrQ57v60jCDHE5Tph3j31jr3VBsw3WorfJK0cySdXVZuhBJHf
lJ7yCS+wBiX7Z6d0Ki5NLlA0xebBZiMSygyHhjADsisEw7bNJxiY1UVSeDh1
0mUGi5i0OQ45p60d4QaY1KRrVhuPNszQRqRuctd9Yb9b/tk8w/1mGvpABOWM
2PHNkfMgOxBS3qrAnCvmEvB8rxK1+vOsSz7uS+cjoUmIch6qAFe4vJxeXdtK
mqI8TakS8aJKQkK9qg3WanqNGNiDdo+PZPGRNIajeA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XBVlevSZnFQ/JQKR3MSuN7K+JYgHdQs21GXQlbnNJV9/ygJQKfj61287/wTd
ZDGmlPclCAyA09A4+YMTIAMgIWGB/w1yM+27ItbScoxyRNWVNMNu5IyhB139
8bGdjXkSS5GYLnqKOMPpLpXa6FXzHIvRJ4UVke+AGBmAR1tnRD8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ur8gpG21b6KRydPZ8uxblfD19FKtak2b1UTBOscN79KYTGtdnopHyeanzjaB
X8vjwbRWKL3e1YOH/w/N6zd8DzkofjB2eoZnp93Fy+HtgirH+IDOSchHXDTG
jTnwRve1XaKtxzgfU1yvGswUlWfslGjW78DzWhWeEPCPaiPyKN7IGAC9XWxy
aUXy6tKExx76iucKzq/3WHdSlXbceHQohr+aAYfxct5KRAI54fGUMxxBKOy0
5uwyK7u8xnS++jOCknrKPnGq3qexjFHIcKwt4Z4ZbkqQke+X/ga5duv4Yznh
nfMKyL7btC3n4zIJ9nhVdjm7Y9xZaXKl5n7MUKEBz3GcKda6titN5RWOxd3A
dAa66c0JA7azw1Uq9H5jsL9diWd72n5piOBsdrk+U4XJfQzIaEpC7lJUSYyT
5ewzY/2PBnmosqsKmruuPiwQ0rI8r4Z3egUifAuWXaC2z5w76oP403mMwbip
fkeilZGIX0B0zsMNUdsMGapnkEjC5UdT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iTLhOgG1inmkPDY27wH0fiKiF679OUv13N44Uer4NyFRR28NDmF3jvZXBDcE
fk3pgMnPPXYFjz7gbKDwk/AHm8mnPQFNZOVrRI3VLO56YJCyQCW9SE4l99Sn
OdueVT69AZd05kkYN/PtYHWYQ98qUi9F50eT2fiQsVsuiEEtwv4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dWSWS9TByfhARb4rBekASUNCu66w1kDEY0KJ4eMeDQCCMwsNbR19OhQXezSe
6WpECf4sGLgwpCVZt4gk+F84mW48PtEPWhtjntgd/5FmI+P3Ooexh1O3Fsl8
Zski7z5j0J4TuIeUUmpSFPEC2ZHKC00e7fXkP33QIyULADhpkpY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4960)
`pragma protect data_block
TOPybO48zgfP9jWGs3kg4oXAG6EiriOPbvWK90BpM+rtp/cNLt6eUmriFgLK
IbYr+iGpgcs3JelQnexz2/mQP9Yw03G7wWVTCwonmcjJRwH3Jn+DRv9wROEE
eZzlkpwJaPREF617a4jrspVc5Wy8HQfI7lX63myR4hi5qZjwMddm7OY59aoF
1pP/g1/Is2qGLs3jCWdHGtcvYP6QNFMbWIozq82vaLGz/Kppop9GOI+T4B9p
uSgs1mwo7QO+YjeE5z5t2QMxd8peZnsFqK6HB6rRyxEzjroCmYpZhb+xYtID
+Xgqv7c6lSpzk7I9fxS0QL2K9BRtEwYCoHmPCPguZ2ou15s5nBOIgptDNroH
XW+bV09DMSGT+J3vHhWwHBvmlkBjOygI8QRVTaZ7Oaex/ZHOAwpUnse466bC
Hd1UNfzMgj5jeMeTHCe0kF4jmQ76LNR2D0NkBmn6r9mW1cJLYyiSeXUCGuSz
rJHjPLaHIXH0fAMfd3/MOvRt5MR55QYwfsKiqwUzxmKUaJvHw3rD79Y2TbQU
2CRUvhdQ5qeDO5Am3JJfUhH4DrG8FzYZXSGQDkAznjglpdCjd6ZSXx/iAQGp
upfJ+5v4Thcp2JcwffTE4XyTRAiizRDfq8FS+t1lerXCoJcsQ95IJXMnNEZp
DEF2etLxF8nig1XtDu1bMxqjIzfN5EgqWsXfd1Cf52a0uWNAc/GHW59L+ALk
uND0DIk/aBvGRtyb55my2KMMu3Wqa1WIdX48p9u1qJJzPQJUinXKDoNi+bkW
hi1CxK9oXqtMilB3qtNWSUyD8xQYUAwJgzM8GgpMGUmxX5fuFmvRNDIZQEU0
FuFF+isWLG/7AyzRZ6Str2EQLfj4h19ohwAPFJ86NpoDdrEcCOIcCw+wFqxL
+z17xYz8pAgARRNenI0gdBnD3sMJv9hDoZYX5P9MEJ5ummSDOIPEleXSsQdM
JvosWepegU2YCK+ssR2HouwAVhptAERFsGRBMgxlYoTUgmRB57P3qae/LgpK
whzQf4oUGkFR7IFQTi72ytn1WRpnFTGxZdsnMttdTsGHJ06bpaxnwyrkns+q
uegyRB6HuUJpICseQkTrzHDKK69XcRjebgEt29PhNGGPTYI5OmZxZGAt4Phz
s52zKsckIqLssZOrxTDVTCloDRWieufamg+cb/bcy3CUnV1OWoBqCA2nYMMO
Om7044d4aBswRn5T0OEdVABI7lFAYN6E9FoE9vX/iCEqE4/7uDDCexeGk4fT
zuyeM1lKt+qUR6dBYaYajoDxf97TfhblLlYsWBjnkgUeWHYQuUY+J/7JBIKR
s7a/e5VTaYv3htX+sB+p9EF1Awl+3Z17tskmtfwCHUutHyTMt0kw27zIUILF
Hu7fgRf3D+9y3agdXXAWeuu0VIgbBzwNINCVApgwJGno68xyDnTCZvPOkyP8
dYRVmA7ojI2cC8NzpcWfieNS04BnCZ2LTf6oskIZng2yKk+RCJmff2WHXMCJ
+g17FJ1sd+0fydW0mlf8u8kWkr3DhTYTNwuTailxKam3ge0wnMa6Laaxl1d6
kLUdPJiwQa4Y3c0EkuYvSIPY1KWxxbmbxNJS7Hhlwo7LEnsM21Lq7M2g7iRF
qUrrCkZEGtMklSj32sbLlwESbXiQ+E/9IJ2ZVmzMEnAX7Kz3JoAKnx+5p1NW
o/M0oX2MC3D3OJM3ku+spAaNrG97Lwvq8QXcc1jJOgSPVu0kmEjScYAa6dcV
tCdiW1sOtw/HucVGA0Fq6tQot4qpZcaAJ9fsSFAPK1Dt6G3v9l5Bz28jHdhf
quO1Wit3RbXIdkatHxtIqXWIXEVOpdgQHVm+c6XRrn0e+Mt2XmTMOFCzemu/
2UKAYNwg2ZNa9t5Fijq56PLOvd/7OXetJXYre+vPnnAy+GWYuY4dX/mkCZmz
AlREjCf9nnZ5/OPMRk9DJBTGkx+UPXzYDKUqHczfDzdyMgSIbsPBLHv0mvpR
jFoA9LJdCUptJR51/wZ3Y9Dh440xX36+B10mgZ+Ck6vT9q7juDs6OK2sZgIb
BQAbHHu4XHLMCzgoiqXALTjNevGIjMtL1XTRCa3pNQUqgL6wFZpXJ623t1po
vzwWS0NHw0tuxlRoG273P358Bg+6YwPhgbrI/G/hsEVGM24LhCyzecokxw4z
SNaM4KN5vlMuG6gj6fyTFOZ/KSB6Owg9tglFOmCFhpTCkEV7US3pl7QcKTll
2kFwz2nbmeEcvm7uiqKv97aIiDQt2oA0H0YHRSzmyb4gxD+dqXVwgWu8iQVx
HGemDgBJpomtZV+aowIJZPowByHVASnIIhRPsfsw7bFfx0YYaaEMXDsW69cb
8jxbohZZHPeU44x4XtiC35hjVVsjQ/3FZOUVlmAJR+YEC/thH1qwEjXSwIof
Pa1CGF4VgTVQ3wR80PIWcsBTLwOhzUdEaZU8eCe0WYIUpZWNiVtdrDp2ixvs
bqzxOomYKu7aSoTpEioTCMh17a4xvsA3OHhtJkzCN7Cjw50DA5S35yv0GCqh
1zPWas4FdXJKh2L4noDmpzPnzdEJxGptB4CVHOpNR4XMTKislJdWLiScPoVd
hj/KYt/5QZZCKjVfo+98yo6/H1Q7VLOs7jWgAuNJJih9K9udhSxebxgSoXYr
qo1jXAFh1Lgh9qy23eIRdBpTwztgCwLIjmtnd10mUYKQncDjGbDHGCIVh0HW
Sf/Sf/mY/gUIRMD6R7raXh7kI9RTGH21g681rTr4e51ykTQVjkzuHeWZQRjK
aCBrcXTPnIUs/aoC16II1/aLlfGJS5MsxCYLoPB63YF6/bBuRgz1JRsysc5v
0E0oSIDyAWglQ8F3TQZDG8rwFKBi8kENNW1LEHkrjYIeKc8yiwviqSBcbB+z
1IWxh4+IpsbKewmM3ERMYjhbE5Dyb0Ff0kusKv13TKCLRJjkDP7tWtyqNZN5
QthvJ+VGXS9hrJUilD/uMLNGUn+zWNmWa9b3u6fEDOrOo3skNBj+Q/Jbp5Oz
uVCX6BV3EXdWfPstxL/zrkXt5+VrHeB5tQuWunJXYLgzfrhMXo+2v8oZbeiv
EUfGaDv77sch4u0NLcqZx06OHA2w53lr0mGKvhS9Gn/Y9aa1zad+OHrNxlhv
FutRUiI5Rnb3joeFCE6gP2dRsSEQxC6/jek2JZO9ZGQiFQdUrsM4zqqb4Eyk
joxPwNtU2cLxQSa4szkAcGOYtxSMCoQs6Ps6507RD7XmbeAJsd0seNuv++53
Rhy4sD5KyHOa53p3GbpmYSurA+uMLc+eIxt54veD482XTOTUkZozM4v8HJbI
YxwiT/+baHAfnpZML0a6xtbW15EuWwi4tdBxvIH7e11HU6buJ9mXxXYRFYWa
KkmBhb3Tpaw7vsvIIWSMEFpJ6NX63DqrFiEOLORHOR5vGsu0vFq06pRwmTss
AtI6UmzOduPyrp9KSnzinJ6gs5HPFc2VpJ1542BFVk55bHBhjW0Ckt1ugwzC
dHFeE74ozZCcMCwqqBqq5XdHtVoXzKRk7ZYqzabUCWt54xL9OVVEZpSrmizG
nk4M8pUxyAcaJ7abJ8ZXEk+5xEkHihj3WulSbraEugDIQwWHZwf49/6xA3bw
4HStQ90xnBHyq2SklqQzzI9wCrAz8mJRlrTVthfLtKBafDXM4ZVyuTMcUeFI
+4vbjXuLypfFEqWKauJZqS8uHwiE6M/jOn/05KZKN+uSUhuGh62U4J9DnZ0r
G6WxovMMNCRrB5sRM2jeFPSIjEmRSBXrfAojkyx13YXqyjBCpfrOnKSxEvSL
gaM4yk9S8HL4YvcWNDh2Ur3sM/VSqhHEob17hUEaTZv6joavZqGJqjdqRxlD
DC8ozCVM8Bi6n3gjZ3MNfj6U9m/s2fCrCP+h+ccF8QuJZOSta+VC97h9pRUZ
jREV/guWhAJO2jCLoB8EiYa5wgOnS1PMEm2l7xjY6zbAZI/uYtu9TEKHQ+z6
BVOrVCae+lJ5I3mqlvo9DETgmYCyL5rfk9Nzd+0+dZoXjRVSYPUFyvIyECCe
O+2ZNn/3wsBcmum9kk1VHRF09XbnNVzTYGZBR8AMAChK17YmwVevrcBEUwZX
GUWpOzbUwPWMEri2ZqakZS9JhbDKp6/j1sTEnzMAyYVoLK5dvHOHHqRYtMQ7
jFRWBfHzhbS2cLCdU+5HaxTtt/z+5LmbWD3I6u1+oFq50v/umoLekOuhNuBz
DVI/AteM1vwHx4k9otID52+gNjZgeWQyKHhwiVFvB/qmJj2qZUmggmhgM4+f
KAiZKNyzPBTVA9m9tFWblmQtQbNQhg68uEwKzJ5LPUemvmXlz9c9mJp5deXC
kWpkNF87K9AbBfaGqnOzm8cSkvrX3pBH01Lgd+gJKVN6PF51S+OT8IhyvJeY
MdxnqNF0TBdYxJLyIYoOtr2BTXsgJpY9rclvgr7q2+UHG5Y8rRiQHSjCUTkX
jwLokizcJ2xXslXNPbP6ado8G0RpxZ5ieLLrlD3SyU/hsos0MMfPNnYNQkm0
wGnaSqOFKJsYlgJgClJrn5FgxApzF01MAdP8mBYd+LiKqEYznp4tcq0aAi/g
VAbau43y2HdQKp846T4I292BMIdFnzB0XyPmAVb8FsZKZhk1GD8yioiwkLMt
WIQsJt7genISMtcr/lfAElp2SrGR9FHZu+giyQv/mZEIPVDQgwFkWH/boztU
CbSw1Yrr99Vq07wRMxUmskuDFM2Mhfd30Njk3ybCvTbb/0MHOcEUZA/byCNM
btosncImTJqVd2ycGJ5SOvZs93Pf1BAdkH1sySgtqFbma1+NGvoW0/3wJGzA
br7R/2Jt5qTVUS8ML8oP8/AKmDdew4I0wG7bJv8fqBTgfq8x0pIq/QQxNvYi
FaWTbRUZod2CKMeCZ2yZJsmnn3HHhztYKDSJnI0xEauq8ThOw3VcnbT1aBRO
cXQrKTmHm0OISUVXJ0SMwfL9dhAdjsieY1OSOUiIy3unhHNAaOTE5WzKE1MQ
ecGtydsMP7USdomsggXcDwSWHESPUQcrsn2rcuZ+25zq21oPMMeTimZr1G28
G3fX61QS0DsVzVTvu1keDXx5kbMrn71aKCW6Lw6IUslN2Kgn4nm6X4UjYbOf
y+YXPsIZ6P2/La1Ev0CQh1RUAwBKaEQGlLNAmajOVP/QyaUj0jHpAMlL8QWW
z5yVMBaEXuS2ZNLH+qL6IlnpXMeTZ/Aa8X3BS5T+5KcDZJTTRw757QnuYZUG
5ZqkuTZyOVN9zheg1qwMcZHFBcEETP05DsADqmFRMN8xF61gKaoOt4+Lo+ri
InWOhr0JXivicoZ6MIsmND+gkhtqSmmfFXGl0IEu78ABliOIsgSrXzrqgVpA
qdaN4dM2VhvaUFhDhAuspeE8renXyQxrbk3ovlUoZAfNPxb8rfukFZgh+dcQ
zsY58sKuY4ahaoC4elrRS2If3qXAtv5Ilu0zVaIqSmSSulrApmzvSlMIOwJI
hIjRI4SunE6lj2pWYVWmbO7yGrXJDyAHUkQ1UBjowBZqU1mrEmTBIE4aMtyu
zOfuOYq0VfBgOYRJYSgPNKBwdetngmPBHHHIUedytj2pttrAjmKxLKePJeJM
u6qzL2eg3bxhKgcuq1pp1zpfw5Xii8mtwh0HAmVUCUYDO9GZbQUVT27GIxD8
vqlP+19OPfFO6ube5dJA629W5epXZV9bnISVis+Y/A35d+KStdt4uwNdrZXZ
N6JtGQ+fMesIYCqrnY3hDA3y8GPR0T1Xlh8IAVgjlbGEM/WmhMBsObB0Ec2b
NJ+F4xoNVqjta4ZOknPlj3xIWeM8SJuBs2hPmmW8Bu2qS5xWUaJAAf969iSz
AoP1DJwueYu0dmYX46n98ianHglbh1YjAwWmxqwSWna29nih939RV3IWXExV
xWXsqVAjbzh0QIBydDTA3ewG9zcJ8kYWx6OpNnlEaNVtr48wWFF9gfPSDVH1
Fyde+BPl8AaSS/yss69ZTLAmVFWGyB1xyDnzl8f41lidAtm2IIzTvlmGLRqE
O5+w3JYkHSZvw/vBDi4BbynCmVwT8Ex4dtlyAxcXL7twTeh5ul863Z2mNVW4
3xOlVHl6W/BrMtYMTfl3d0NqLYQrjMzK/lz46HD1u34Q1X5kR8RGPclGddPH
XxJhL1bEOL8QeoWFf8X1aUhtmH9Kzy6NlcpX2hYVNizg4Bfkn6TJytSH4kQn
RAaF/Kbu+xuqb6y9QItvAfqdTHsmK7+Q1eSy7cgOsGPLWZC7UzxbIPztr/QD
mDRQcQrhcMDl/jfVuqWEjQVG66qjQDCZpmsoj+JkHVgwvJ5afC/qx/byEW7S
HkT5dQD+Rk7Bw+jsSh87UTJ4M2hj9KT+hobQgGKy66Snjlj6uUkeDcle1Ni7
Uw9U27SPt1vi9cF65JMovHD3gVPlaEj23HlkwnTgP1W+tNFBCvL8BETiBhFs
PkJjAq9swwH3ncwI86ZrWltn2FOAalojuqkLhiste8Hpg557/Nh0q74w1i7/
V+WiYE5D2mOyHA42wRWLmT1xUDcmQfPYg454ynacw7zu3gsaJUefj5/Vno9g
Qg9FraDQzpmcZz5msukpyot9F23ZHDCFYFOJWAjR/pXXlyfr4aPOoTwlNRA8
NIbAh0OGMdgH5A==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI1iFd0y8CaFmZvuH4trHLDzB8FWhoKyv/eVWxDCRT9GsZ4O69ici9kevwDAuLKVr/yt1Q45RWMh6Cnme5iCvTuqDo2Hw2bpT4IVfV+onG1kf4vq1DLN0H9Zz5N/NNyq0k7ew8Y6fW85zz7TejMhWDE+zTRu45EYCzVEcIfdHclBjgQlmoBvWFrCbbC/F7Xf+hN54TVKAnZ0BMwBIIKQ5c+RmFd6/sM4RKvlO9t9+MBDeZG4PscIqQ1Ct2lHkinlFUh1BucdpPS2Hkwt8Eak2ZvCXVasNlGBxc0fFyhWSNc0um0G/hwgRHn3cY4/1M9g5meudaM/XNb7IkF7olf3W9ru7fJ2GNyh8Ij3TMXtLuICDr04/qMdRI23cacod+dvZWF+IpuRaoZW0tW4fUJQ04j5FCKK/WRlS4qwXJEywpT0vM9Z3gilB76vb+/Pnq6kXIMzOne7hBsljWw0xSACE2WD8d3b2ePvRfqA2vEkwmySW5IJUw679oAWt3zdD2oD9Jjc6bmomUaCnibOe2o7r6+kpwSauE5MeKjfL2/t3lqzZARSZU7TjbHAWh9WY0SLP0ibFdZfe8wJ2lz6iEXgsmNfWQOyQga5w8a0G35SlfGI3hADJHyREZFv3obq9PESIREffJzQ2qWqefT4Hmc6i+ETl3d/bznvsGv4QApNopkNyT8GztwSSPYh91aQIldF6u9roa+O/9+IZiYtUhUcZy59qLn0Gysh/Onq4ZIDUDdnYab6xYjDh2ioio0S48Y1AqQCuPasnh8b2t6/hz3vytaS"
`endif
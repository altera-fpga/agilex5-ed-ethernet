//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sgbVDPtOgvvrdzR2V64d0YuK1eZsBgZx8shBbSklzm2axAPUSbUkr6+6l7e3
M+FKxUgCQ2cd87O6/JDgbLXCKL0hgRoicVXIs6CwPZ4gpwWfMSYoKgjnFfnk
+1HgNaK8HHn7MgINthtX1w9pNUIZR79TL8rwwzZpbceERJwS58dbkxtEzFM1
8gOS8devX74CIml7HmBnpjzaZIo8vQmDoOQP77xOkuOOPn4rWgGN/49MzjAv
66N8vbojq+AnrUH3FFZxGT0whxJbQ5G/JHRUjNKokvIjO9SDzf4kn+b4qUnd
iWhzDemm5Xeh99Txxft9D/SCa39+yNMpO991z1gU+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eDRkqsXjjfdq29r/+WM1G3RjERFpQLeaPe7vXUeL5FH9Bsq3467BeymM+67R
O3HOlMzuGIbLgQo2Obn9LrepOB/GdASLPKLoT8iG29zWrh+4IgmgQwDMOpF/
lTOtnxcPvYsWS//Uf/xSqDectO1HsC92isXXlU3pPjibWIs/06pi4hWiaBJD
/nNnpVhGwjuSAWICfNR8shcyX8OxIWcm7c3hgRA4YjhrOt26mToKcvAkEDhC
wdY/MS4mVYUvkBa/xfQcsygV4WGmRYUquKznYJPHPdsoPvCzLkvRofnPmEv2
1A8OOEsI2ISVANn6ahik9i4BiyYq/YiHnZn3jYTidg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EiscOYOxP1O7WMtU6kOa7jvzboJXCI5zWAgwchuZ3jurTQLvyzm5f2hP8MpL
ruf/BegRw5shcaPw/QRpM+dwu0jilgzHR64dKFyHZmogx3P7OSXqQPzZlFZZ
43MqoeSgc5DomCI+KHuOls9qrUxmNgyxbWzaMsVHZhRpsH+OrJTvUCLWOq1X
vYc33r0OuWcZVEPY2tifcBQoQPQDTzwqUT6xg4ycr5yy/81bABx5KKJ7oFfe
x1GMVl4L5ffvVwGeRlBmpt6S/n+XsBpSQ7rHp5RDQuxqe3E1w2GEKCoXX3hj
c77sliBCUAVCtFL7pigVaDCVKpMCh0VoI6ICoyyYtg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kzyai8cZcf+JZ9sllxfChuy3WwI+9WICpC9kG/r63bCRrTQi9ILqAhgpiPTY
4sMFdZBM6hHi9jHe0Pbm99kGk/e1V2kJHTKXH10BEUhSee0e420BcvasWJ8K
xVWHdpKPGfcaB0PtYadtuxdXuvgSqBI3mwDOl2P/7iernhfiIe/dw0YOlhM6
Ds5GiQw1tEz/dH2Q3SAP/j3xYXu/OF/fuO0o709m2u3bC60NRGKilaIhZ55j
i1cX+Rk22H5X4YgUlRR1YcMbRLYjX996sjTxG2N7XgYUcymvHSROEnZCmlZm
T1SQv+zfthPlz0hsmaq+Y5vwokOzocSm1zrv51+ydA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G3f8QKV3iNnEZXe8erXSKbTsQmSFiE6mBZRYVpO9Tw9eZk0KNDynrSok2dt+
sXT5469vSCSdgCIZNHYPzKPzWw9l35N18om96ipr+Nf1WuX8FXkHcli5O/dj
7ZlCLRTtMt4WaqO++ao2kxaPnQ4PCgazr6C0S1YKiEf+S3iYU/g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Ae1+jb21Yt4187+/TN2kks5oIKqIcGrqdS13FxAwkbS1UfDUB1/8too31N6d
oeEzvN3auN+kkyk9Mq3VtRuOsJS8K1XDNvsrsAUBHUjLqTAxEWbH1rOfJu2z
IC4mosC6GMVDwDSN8ePBOiUVZMjgCSWKXk8UpMck4TEn1J1ts3hP4b2qlpdc
R6efyVuoUfVfkGbkhNk5hg/dILSesbvbVPokE3uGGGcrcGoL1fbL6UokWFcT
utCL1rqL/0DsnLyHjd2u0D+8mQ5PUu1huq34pzvlTk9Y0SJeT4jPLVBLhxSn
xz7Z0e071zkIFTixrQ1EiaeLdoWJA78iPDzQl6SdeRwTZLza2FyoDt1Kd9kL
p28tYLawKb4E9acbNNAPV61WKzNMSPzFfiSXMNlkASYRmYIvfuGDbI33jDZG
qmn4pnxeWf+xIS+OjHwVThVZ2vJWoDKBp2IZZhRaVlgtBkiaAvA/F3IyZd9K
osklUvqejZ58isnaDe/flWprpSRx65kX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KBXwqZJrg8iO1Q2I05KM5ZdN5KQmc1SsWQvi68hV3XPKqKJkPOSdLYwHHjZ4
w2+kVAnDlg1U6Duap+ga82kQSz0xrWFs5FnM5j/6PK3iHFzZcAzFd3InCrfZ
cCikNvW0hcxzO2tHpOktnaJsZtSBRk4bT2AbhRPouHUZGVKidSQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rqnZraXj8fRCBOgI02vJELJ/pBSGFr20DTMfiesRGu8mGnBwSJFY3zpeGLDN
70mPmJ24bVI6hie3EIMoLkZTY9wzuVwQ2M60SLytGo4bgnYV2wP8YvX2ccYp
EbEejTZgkr2fvRtYF3n9bIiJ8MFz06m9QKnkfPU54ag51dHKWr0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 64464)
`pragma protect data_block
+QK8uWjqQmXxYAQkGU4KGGDHmwrdKTvJzDa50c9ssAlkmh9yOiv3aOpXPD8Z
XcmrFfRMaIFF2h+qehkf0foCpvuVG3pnfKeIJqTE9mN82o//y9eVzz4MkJaU
k8+/xSqVty7l660N2nibksY1EkX7ZDoWYXq0hD6EtVn5XpRPZxr4G91HD6JM
GTeIGsOa17WyyHm6czYSiD+gWSEiIMxWfNfCG4f5OwXWNvKJAyTHSJP4W6CG
AAMeMhjcqDoiKyeChvPFBIXhE0I6n7S3PY2n9iU8De7gfGKIgIKpdAP9bRVU
5YkJqFDGowFGgeb4qaHHr6ZrsM7xnzBDaGRlB1DcuNKHfYPVDA0OS384xoT+
gOvOBOh6/3iVQMJH/JmVhEhE3L6v0iB0e08pWWPzUqcDB8IXZB6B8YLDgVo7
v1n6HsRgX6WPkC/zdTInkoJm1dwhvx2/uOIueyB6e+YT6TXIuK6X8d27egCu
7oqR6UNuv163YP2klUvD/r0ZHUR5dAy4L8hgXFf1N4M0Zw5gF3IDGVX/dBxJ
amuGEZZkCSayuAjIeAjL8z9wcRUaZAgt9pjtJDPq+Lg8PhPUMwmzsi4fSPFf
hpxjSQ2cjhMiK/GLpKf3hLGz6hNhUYs4dTtCSyZlZ/ZARLKIsiusT0gobUMh
By0q6JwS7/p39LakxJYWSD/yzV+dXqb3cf0+914qJFta//4ysgoAGxSggAR9
+8e4YRBREv2/CUFBst9DgFgE2gE1shFji9Z2e8JCNl7wDcWoYU5IPkQCtWtP
N9rH/XWjAgeLgkF9R/cUqEW3y55x1/zAqieYO1+HBuefmDb4MIxvLULGq3bA
umkJQeh6fcuqIrsU65WGpwPXd77pCmkGaXohOh5NKEA7+JUYD9yDKsBMSi1a
xdBBhJxYDtUAN4rnBRnAWgQo8oXAmlXi2JTuuj336Q5qTYfI02fwWP/HKgTI
lTVrgRNFRm3GoVYwukjtb1tguDA8GcYM1uk3CVAXqlGv13I/I9596raXcXmW
jquTI5jQCQBbWchC8CMiHcUMeaij4qzwpslDI2XCtMAvMgqthDiiARyvF1s4
FrcTZFPxdRsfdSqYGuCW6qSd63Nb/MIVTBKJrkvIh+SYEbwBRqXZjGCONIkR
cDVleDLmWWE2oZSpEHC8f3ZLiJQEwwPnToXESCqQdwEXwmOtUh+5sazkrasT
x7+Tbo03vgzipDJ7j6xKcs2EqLkXgVCXS+fN5ig2VO7YQiYTmeYySJ5ne/tY
AWzLbHlJIAqKpk1t3XmNqqVytMMYNBbTKmlZ0wglxm9+QWUgMy5FT0OGN1+t
RsFGSILsyB63wklNmQw50mfdee5+KboF2P1olNycZE4KOGE6FIovM77BWlTY
Mw+Ta0Qs4pl1Bf0/8+Ppn7nWCiwl+Bnz3Aguu00iKXW8SGa5ekDpJPFPbraB
X36SgtVGA/hzrreg1thliTRnZI1W0lIFhAhmQnc+U5qhaco9c6vi88q7Gc8R
tzgQQFsckD0UGKcIlcxSfRQ0y5Eq/8hLaFGEt9JuQepCgREU5SJ/64frYclO
Ui02o4s2hvjc1740POBHU/u4EqSuimtoHLxQxEfRri2XvsaXRDHVd+izk1Zh
adj3FFcEvCiPx4S3eTBZn4MtmotKDW/qF+tOUD6bc9w/ZG6BZ49dPkkmmrkv
yjncV9ni5oXrEeEjh+wboZ3KP0RpEEJOqBBYclaAfjYfIKPAg/DIsD7X5lbU
QsjxLiHvHAO6d7bDW6vX1vDhCckV83GJd9nVd5xQm6DLOQhSDTHbaOSO4iy8
F/d7sBYptYse/3j/WGNCOLyodTAt+gAfDt9LkUkreHu1Vp9btgyzUQ6qyaSm
41MLBnAXc2PmSjs9KJevTYLMwkKIe49DsI/racgI9ff/Svs0hD2RfVo50+fd
oJZy2TRL1iCif8K5raEL8z+8dA8hT7P96peWFVDTbaZkfQe8HkcWgltE7gkc
JMlXwu1UnJlav4mUNTNmLpMj20V9yRdT9O5VVjrd1qFy8cpY3gIVbXPCqKN5
GqKaveylSwBHl7A4ElbZdyL6fcb6S/21wAc2JpevDZUymTNSPpluhQgzl0jR
xIxUWKFNGIBGwfFV6Br9920Wq/EUTxGjROU0+ek9b/RxyXKxRF63fRCa0moq
YEFPxjwouIEMtgW/C/rYfNU5oayJiM7pjnpffpoudhqs7NYrHFmbxzJI51s1
1ADuHuMk6q4PZHMbiFQuQ+EIv1dB5w/mg6Xyx5SYmkmTkhOebkOo2IvqQe2m
WNJoF7iKHLNDWvBn6RKJlcjCsY2CpWm9EEiY+fnWGVJQ/8WBIe1q3eVlMNTF
HCLjJPJp6AipkOdThfNmiQNE7BftGIR7GdaCDhOG1oKtH8LrcYlDqWplS4Ah
xjdgTUqMCVgBKzgFbP1aBMD1N4Hhu57425pUy3sNKLjGFUUXeazN6IyW8A1s
5ahnCLBT/FoeE4EB/rbupD+tg1uJ/h7flskup0wlJys0BBqiQJ2Ox46/ITcs
o1Esina21DxU+HPV37IFv884GkfjkFcjF9tlAcZbEYgl/A5wTI88ZamWArTz
TubX3poRuI4z8heqDF+xiQ0UUMjBtb+hMyVLLVymrw+zqdyFC0ija4CwPgGf
wtX4Gp7G948Adw2PJotxghSzMuiQWECKr7DCR8FGNGehKl8i8ffiwheZb93g
WIcKDKq1xuIXf2HMO+lChDcQjqCCFfabjrO1PBOj/re6YGHGIHRgtyBiDKwl
meRNZ0fZIqYaYTV7WEATxIai9OCK5zNRUb/a4kpXdBsL4xFYulNhyb/XXFuq
V/oET142IBctMHY4ONh84yDSMgYGDeouKEIr44McIQMeqF3koEicr+LdM+Jg
LJQ9Ep0BqPYB1nu2wAM+iMXQsafvOvPsYYdR+u+HVlZqUEOv6i8W39lfo7zA
X8qgjtwtWySM6zMoQohFyCwODJQ+Unsvn0Ev116zuMz56znqEJpA52uLnaXb
Bl+qE+s6Ir0g004EdDw8NcC4i+95gINHQUwLEcAtY+0/X940o8MoMsMKWxK1
SWYblPMAmx9H7rLEb/4kJBPmlU8/axFtAnTFk1D0xOU3FVg2RzUoiJJhI84Y
4fS4Y+MRqh6+RzlDjigrvsZhPyW7TG/vyNLylIHpj5Mw9+4H3RU60xuWjNty
3Ll/YUw1J4JGlNM2RhW9Uh0dZx/Jc0z0XHSIBaqHpPmh4wFbcXWVg/XKzU0I
Pg4w/QubGyhT500bFwIBg1nk7jBz2zr4Wf8f9JdfqIvfUf5MPSHgiiez3JK7
xSyqJgIWn1t5g9gZjHOThI++F4taHcB6fVTHXnKeI/sLLeyGdOVyVSBBiPmk
Bs21SfyLrOUSkkBBBZldphNJf+cOh21DQeJ2aLQscIaNIHHn60bNKmOuf3pw
EKd3nAH51o3zOTwdqIpywOz7kWUwZGPlsvHTUSIrLv4D6K/yPkhqacNaURgn
EaLHufNvNC7Crru2jiB5QAPccyXiK9mTSIFDlisPgySvERQfG5/7i57sb4C5
rFyOluebdeD4X7zo3sr1DOD0BhsurRm27P/K14IjmXmER7VylsnuG6vNNfWa
SKr9skMLH7nOTTaOZy7UDXBT3Z0hdfD53l/EC+cKQ5Y7HowwTe07Ag3m9py3
jB76swZOrDbWX2JfVMT1nZJer7RYjKCSTwX+nfydhCgF6FrMLw1tG5oXBVVk
FvzptjUEpbgQsmsDH5eskANu9iHSIixZ5+s1ZitIe7kvceYDbphxxXCzE6y+
4ptNxOhm5OO+BH3grALfVvZQ2Bfid7ba5jNEnVVlK9ataefMsKmG7T6enWWQ
mwqgns4nWwQXaq6rUvuCHpyCfJMdNkNqCG3j5FzmL3PqCdjJ3gngdZS3I/wQ
NYDgcuNNYjoFqdTxsNF+dp/XTZWu9IUu7fbzX40Liy7o3zT/UvX5r2116vcx
BJ+rv0VgzMaEMnwpoBlIvXTGWeSHbhhV5pD8IBaoF4RqN+x304Luxamy5bmZ
68i9S7enrCjr0h3w2rZwtabk6IsNOQNqQ78/4BxcsE7dm/hRAgdGmqVc6MMx
oGzr7s0IxilkLiYc0QLhDUZGKzkTG/Tgqhxlvj5EJY0W5dVKD6/79/q98Mor
URmBd/6ZmFPURpf5U9Zgy+sX/qJbsPSQiAwE2qymbtx+HJ74+iUa8y0BdJuL
NMIvhmM3tBi5vvxa7XQl08RRJnI5+GVTMjvtS4RID5ovUPi12VPj12fyQNYK
4Qu1gC+xRITJtKU05F9blALat5cOQKM0s3Ohy6vF7hX/xYTsDTweRNdPwn9i
Ln6OXioT/ysV8eP40diR0FMGRJ4KjI4Y1dirFmZGJr+oOsC4aNLQr8QlQyqO
AOwOABLla5/8TD+Rl0w17ZDX2R/tuoIooPE/jSNwfCMUcJfBIee6jrm6Aohg
fgo6/AlTzU979T/4A9MBx9gTKD6Ak40PjJ8WrXdDqoXq4OB9xsdzIraIwk5c
o+VeLboz7lgOGwZDvTTd1plbOL0noKYoabjBGsYZ97ulqyFIK253nAbRGq5s
Q29b1dZ8N3iUduDchT7gbBHvW6fIcAm7qnYCQ4gTqs9Y+yTJog2HeoVhgD9U
6OfL/lUkM2mvSEH1NeLLXueI0Hxp1zQ3VOaNQD5vpATDDF/h5sAcnxL5orbD
EOcogqAvO/WPOP9bCV6KSzfvlJoRcMqqsThBlLpvXxJKVDqaZYz9vho6cLBz
15ApubJJq5fO71MGNYxmLZb9Q7PmUAyaYUG/IJ/Br63WTuNxzFcKm7uwiaze
RQqMDdGy4oueCQeKdYaj0GUp7c1jWLXfXK4TtdhNlgJ14bPxS7XecBHI1fAk
TFW3PeMOmraEDiGadLd5252fxXBG11eXt9LGM/pVABn4/vIrpwVBtY1d5Xue
MV+R4PqzQfHisL2TQd20LZpLtKBwIlhyOcP766nyS307vDVawEyn0HUCoGOl
yAc6wfZcMR4YCyA88GzmlYj4/YfGN9vqFzHSnhEjAyHTq82QkOCIB2R6rU8e
T8ZOU6GLZ4LHmOdgi9XYA1izuqzfy4Ve1TMEPU32Zk+Z3m3XL/QcYFu6O78h
7mttaqpMfRXVA1LhkoamIsBCfZV6P/IlWQq0DtnUbU5hz45CjCivgEyTm6Oa
Vle0es72E3LjLRzrl2/oOIHNue10JTxXVtiWXz1rsqSdwGGePfcVZ1mHI/l9
YKQw8BH9UznCxtuLnjvHgbzdrkoOaDeH5b3EzHDPCrgUjl29Nu9Ma/ySEjL5
4nKTjypD1mD1EU/D0Zt2JUFwfzp/H7lwKPG80J0VFskhSLuz2Y7E6CiNCrQs
FzwPtuOIUzeK11DQKrzt0c6AiCoe82SxX8kL8gyYzAuR7j9o/EurTdR/rTUE
hiICnUIKBeHc89DuRMdSk297IQub3mq0BlsrkLJtZLfmD8UJmBNhww9UKh6P
6UMBknD3hf/L8rFRyWZ8D2Pzvm0ePlRIKaw5Gytmv7Csp1PpaaRYOYR+JyU8
wf1oeeyoWqqgIswogO5EBDwLgeUn/Z4EdF95Lewri6sl0yAym/mfwWkY4orx
ppLQwbimfpkATqJGnvdNbCQ9kF4DugOrCqGCeqTzfkkLJHpfGF/s4IESGZCR
fHCuunPuvEcRnZ4pfn2TjE1vfSnbPxPdeygh2EnQdVs2CWur1uKULtV90Quj
CV7vBn2LfReXCp29XSQgy20NxDSmzFr3/q2WbfcSB3uNgJ4EvHK8C6rToVGe
zP8hLGozVycyx+Ilao/5/SDP97yVoo5TT9BCt7hhbFlrYcSlTAIouhzkc0yI
RGZla4DPLJVKagX1mddbD1xP8KW1oxJtx0nEe0GZcYW5JwxSV393PxAMviWn
Kh/4+k1vJQ3PUsvboeN5J4XIXv5KClWI4+UzSh3KMLLz0Pguhnw6j20/APbw
ql7nGDjwfISTEHvomrOTvSWHV065yQOSUlK5Js4YjUzdu/YPLx2WJaTGWxgg
V/PMwFhzVzL7RMqBeKUhH7h9TiUG85ygM2VLixX6LatZtaoQFILfoWvXjak3
vcCht3ZoWY/qhnmKGje5blEZ85+bfBUpNyn2LGpbTt/t4EZP+CqccaJ1EbFa
XjdQrFLKNhO1p9toB3wnzEdtpr/t1FukrdK3jgjXP4ZQ1BZUR9q0ia7N6bgF
yC3zoZndzf6V575G1LmoIzBqL5x+1gf3v9kM2ktgcANRhel45sDn9u8rF02M
dixvlr2UCgEvRkcAohcFVdycnS1V9+r/BJrpyEbC/C/IUBd9nR1V0mxC4JmT
jze+FOrjfOl4mTRGDL5IhKd4KmrBlqwmqNUt66UxXqmusVn48DRTLdcb3LZC
V++7sCdoAsgfEYGeHaovZC+3FhmoO7EcItMZ+HQi4aLFk2KFsqHWA1a9yqOR
JkA8rzU/k0EdQHqLpPw/xD/p5/SpO5uGd9TgV4uFOs0C9BTOwJmRCYz2hr16
GJdUed8wK0nkAzS0h9OyOFDdWAUggI0VlnMefgsQbQsEoc4vpZRMR8DaZJIx
oQrsn6Sqi/4Z4mQVvQ1HIrmO0a4pxFZLAvQM4Kg7/4JzMX5WIysQFJKd8Mpn
HdBxYqjbXDl0vRp8mNqiQD/MHiLPGUagc3xcDhuVvcV7KOTwLy5FEu69AJ+n
XgdI0GkGUHFfP2F0389yqc4DhLMXz/23AA3tOyO1jnyqGEYUPcV8Gwyl54lA
gAM6NKa13WyxVWdPT5fS2j9OubIGA0IC9p9OFLa4N5QO6ocAca+FjlfZO8VU
hbNDGsS61rE0WR81YgnyuY+gkuAPBxuUHeuhXTX0hRXV3NH6j6uN7pCLNrb7
+pRxb3UDJO2+E962YGTWdWeowObMfD+fXRqo1lV5ZCnc20ifIzIdCUi61lKL
BljvpFxYsQftHuqVGoUrIYdwXOpZesA9jrympCD24nYVGTRMl3LgU6FM3H/0
4gWFVWMrKfJ8BaYRAK8FZCFEs5R5oiUrTCDv/9kDBDapavCSRvg+Ylzln2Vv
eBsHiAEySnjCao4nUY5rn6AxqRkVOBapwEFVb1MZcWX/Wm/7hOGvqkD32F7+
xUHBkGM2S04QK5lBuz8ZscmrmhJxwqNLzL49s+bdo7mAEh28vxx5uR8BVR1W
NYLBx1lkvrdiHd+BWdzfGKMR+pprfL9arCUykS7XpKAz1WINnu5Q1c+fU5NW
9zDhIesRLyvSYrLP2OaBFXfRKCxPiacvKH14qZXdumChSLcW8NkudiT88zkx
bsmjD/Iklka61PVr5Mhx0eXrovrJTU03jJKyf4K2bTljA1PcebYfx5fycxp2
9cc9twZ0Voz6L3EZdf8osL3sIqWHiCPPi5Mao4Ta68lhTFQUVDdqqMopEdSY
CZtoMfV2jLt47zavGT2mxLKU0c/snnIAbd0ZMLj8cWF3PabcYLFgBWfsRU08
ow6/qMoRRQZsV/ODTog+QRbb89DtVqFTD9VWNbVDmoX6fd9B7QEAPg7hEGEI
x59rD7QHo6FwTdCfh69zIIVQU4cVEHY8JoP2nDUoXoOAa9clLzVZdjvPuJzx
SNa6BnfEqfv/Oq9c1ZKYDCUMgjh6z/wCaYicNefA0A5DUpNslw+EuudRlK3N
wjTx0yiEhwE34gF8OXtmkBBAjjjsm+xs1OTZQEOQBg0HDuaJ6U6gp0HKDfcP
19AhLF0uY9NTdbS8RUwpa3SCmP2vvi9A4D6YQRZJHGb4pm0RwcTHd9z0qHgk
Rk/gd6aFhJZ5oJGV0i2+Q21HaOwL+tVrt4T4ntKd8x2d3Ab2X8cwxh9nwWng
FAWfTMTrPhG3h3LHfmjWXBmbqYHAF7W5vNdxSV46zCIkfmqsWmRQ80GITt70
ryTbSavDZHuFb0tO9nDtVyOaMzb8O1YfW0SIOGHL4BNLfYcs4htZsfD8uFiG
rvCVVxaX+JcdYPR1ldNmIPVmdVHV2eqbWf4gKMF1IIkaoOnirVsSh/JvsLUh
fPtCFvOsuvthX/K+55M0As8kVcAMeOWsqsytKt1rN7ytRaOZMfMh08+o+5Fg
GIRQiQyQdTO/iYGIU9uoAUJSEOZwfKwDAtiSIITHBAQZjEFCn0Ssc3IVD/yg
Bf4+mXkTvXeztC+9UziL2NA9+rvohEdozkqaxYR15BA+wg3kGnvAWR5TnP57
NZh97IkxoCGEY/fK1DNSmIFVOScQIpTRSo5j7BQvxmGwawnG3tCKAvION4iq
1gKJQfdf4CHHNgPAMixdHHsFuIOgonHE9G6lOJ9rmZMNXY53LG8iesDC3pb5
VQmu3KpfXAatVIwwjghYkJ8crDfdNjU9jKecEdVHUzQX4z/EdmK9eIgA8qWO
9JXiLvzqpcwKc7lUlF46hyoe6/u087bO+uFGbZCO9RM8ZXZ6P/eeEjripa0m
9cwzOOxa6qj2KgYUj3Av3Xejt8edjf9aQ0Bwij+DdnXjOZ+ewjLutviHSHm6
QvKWrelucPhbbTyzxrxjWE2O479Tl/1HjyR9GdIjpqEwRyPL/a3+8lRDIBW2
hMBVnW0HpggZeugkCg9kkQrKu91QK2H/FGUAxVQ3k6LnmVh6syP/jwnHs7qp
5vrtA8rZc7ZDXNrP9daydN5azV25buYvTaKFJFPTR7v7wZJdmIertFZhPJuX
JnQhL3ZSDMSgF4psqnO/7ZKg9KWapTnIGeF0Y3Zhn9tqrNrgFmFtvp74SeGs
kbYESUh1bcwtvqRvhqd0Mwf+CdSNdrSD/F1ueZVL/UNKv3aKWfJPk/nJ4RwK
NVzi7FHHscnRPYVpZvtM4h0XEG9zSZawff1701npYIknq2zmQI8sN4fAJOgE
f61XtuGy498XMj/Mu6P6gHytMrI3nd4VIAnkJF7K0JUht4b6xYi8J6LPPZCZ
4B2LBakB3OumTEAKcMtkzTs926t3xhWJq6Dmh5vvbiQ9oB+zPkAnPxVHRioG
0H2iggIK0b1+p1LJ5jqdVVbLHbEDTE/ObnXBMtr43yUM7VYmDkMqoMTr7kpz
YU2BsKk4yQAv045kgBsObq1anEBvhdbNVghBqFX4MNudrLT5GN/eQVWNoH7g
H+gFpVkKd91GXA0gbpP0Z7Y1tFJ7Q6o6iplF+d9khczWNvcjKmCGiU7Q8e5l
RHXL3VHKHnRJBl6TCZXIrT1DiB0lbo3XhvxJ2UTXBjHrvBduAEPJCK7Hbwfb
2nuDYQR97bQ+JgelxmQltFBx0wJFeNvvqS91dU0dA/Y/uieNqf1rCKEbKJaM
gXtZYjU/d2JkHdlrjlAyCnsG0tqjsSQqj5mFmLTDgwDKh+t6wyOhMs1xuCXJ
+5E5qQETxUQaY1n6HTTnv2OSVY9wVhOZVUFjT4JgSXyyMvqXy20ZRe8rCU8a
atYBQ1vd2PlPb54gi5fIwTfNObBPnhKRJcpoCTUAJmsUdzn0XAFyQaodEUBf
gAfrcEzCUklzdTMj21KGNQ70ixb0FueszyAD47YK5qac2FRcZCIqI7HbtEFm
pvz22zbAVnwGaAyCUwwGVCfdJ3mW1lGoxT2TWHyd99gUeoKmhm0DBcbs3WEA
P/ecOma5ZgmC+eZV3D/X23NH1FgA/aJSFIe+3t0UuPMBveStp6fjnwHE15HH
ywP0JdaqAg3ObmcDTUGQWMi/9UsTVdFOH+iLPNaQViuuyOJzHDjdKIePtsKI
3q6TNRqHKbZm6WpO6+iCI83LXKVoYXXVXImfS5fw/cliuelAUQMI1QAaV73K
TrPMTKhZ5j2ywX8YOG8jrynjD+CoWr+GWPN8t7REH/NpkSvYyFfZhn0MSL8V
tPRoIluosoghfz6r6mZjZ1MdrrirFVz/Rmb36uUsWWXPBoDeJD9quZwsrMBb
tbNPKsJQEB2zlm9FexFkEUYBR1qr3kM7gSa360WeWnxQhZciXGw774h3dg8d
5CwdFDVL7TF2o4kBJ703qwxD7BWfZ0eNe279TTt1T4lNdslpaFLWT6RMNQUO
1lzmCih98cmcXaQhIFAA5TTP+hGFaLDMsvFakH7UWVg1BC1hvjdJNVnWCnUg
MneA198RlVmw8VNtVYNFwsietqFvv3amfkMs1no/JgFD3a4K1Wx82FZe8Uk0
CiQBlGEhlHvzzv1cKXZMzXZy+Q67dun2H+uYP0L9rhUjBfUW/qtkQTIzaQq9
j7aaSh4QEknw9cmxU4wj+31n5FVtegAQNXdXLUkdZtD7NZf9QRe3UeSTWQlF
MYTOucwdrpmDbmmTvrGPEb53gigcomKU+b6Kl4U92VfXTUu5uohVeKJ2YyXW
iuehl7zBceGtCkHb/xfSguoK/Zvmcr/youA+Na3xMFH+cgWtiyLyqshBQPE+
bMMPs0sFezIwpcj3Y6q+bfu6FlL7wsf7ehZR9E5QA4sAGt6LmWPRHUzBBOsg
fGWZnZjhWfFYwgC+oguld2f75l/Vm/4PIukcaPvLCmAfm/ob7wvMw/S76IDI
fK8g5Vq8jaYE8G8r6QaqM1qJoFTJjkbpDTsgHJKTgPB7nt6JQeB8d9frlUYB
7k4M3+pkcHQZLAss5AqiSy0cOp3GwTWY3V9RiPJDhaCSQE2VhUXW3jp5BaKN
NhMzmlOrZHCPcDRWeTCwuzmCfXW3hCjVd32BmN57OWQ0+WHImmHt1+fMeq2s
xCgFNXymRfLD7LRdza9dIFvcbJ8Clu+y0Xi5Nz63vRaMwWbkwCh9SXTZwHTz
EuudCJ4WfeNwtPYiwE4BfisqrGg+jpmISawTiub20M+IrT71C7UF3LGhBcZe
Hr4CVi9dDOuiAg9kQ0O2TYwmCAi/nvbhL7jXPR+9BQzNWkLlDPe9vFGS6YSP
LMPbkhpaaR2zlTUnAQwZ6OFUSv1g6jG/f4oq/coI97oHjYPlu4JwhhISJm27
YvW8aXmDIggWoaFry5OIvxSWisQ3M8UlDMMj8b5AGr22WHdzX8o3brtsShST
JO44Q71d1WZUP56DtVmxr2zQwad8i5pGXQvKiR3fYA9xD9Ur5UdO1mIhAuxB
LlSzOGUaVjBi5nocrcCCl6x1u3DeLyMufy9Gv88JlQA9KrxQlU1JokzEfRgi
77pY9+4IWf/U/nyn4MtvC4vnrdM6pYw/HqF8t2xY7xjCM6orIIVEySW0OqJ9
KKKpNx6vTWBNdzlNSptQW+nmx8uUZeqfSNP7I+ckGAMnfzfegefnDnrVWWiJ
/iyxtYTp/s8EuFfJdwmiH/tGeaLMgaEqA1nKiHbCErnsEZUEyXtx3oMMTafU
lMIPfFvDkqEMUzJdVTDtRuOCJkeeVCkYxy2F0t2mqYowsuRlxXNlW0KCJ1cK
o4L45d3sDMRWcsPNfojrIvk17d5vEPRZejgQSsZu+9kxDDLSclUSD8uWwo3s
+EYGBwMy1QINCS+ClJq9HiDtaShwiXVXKBKPYz/mKo7TXicg07VfH/CFzRhX
rithfH5kTYcP9PHkhhlCP/GnOvEBBIK0UsfL6PhNNzI0E8Vkphcnvp5R9IXV
Iw428MYc84chpbQr+d+lSvMgT4gq7S7ItoLzi3PfzQ5xV0roMH6yRC8m3ylN
uasDaFBDCkzbqd823KwKSjjX3ksXAUF79/HbTSdHW3W8r/YHV+YFxcsHMLwI
RwGssSUrZw7ZR9GN0Do0djo1rxi8ppKvo6SDjv5o+a/BJkl24tryoQob1MKP
FQL4D6E5V5Md8iPD4A112TE5sbL1qms8fQd/j5hxUELTzcy6Ne3q1PUelDn8
xNuWH810u2Tn7h6Im+z8J1j77+iohBRiyGrkaY0HXCgEHAl/HtestOKZ/Hz0
BV45f3CLaLnJG6Gi9N97qGuRkWOFwVXApqhHU4dRPV9WXq/sbXeyHu6ryrUs
/SfqANvTo8Lcl5Uk6ZBUyBOkv+2j/ZSv/ZToWRw5prTcgBfNYFd4DwX6uvF5
ois6RehdGlLiUs8QXO9RR50Hcuu4HG/l+wcsI3dS7/OILVIVO5jn0fuSq6T2
AU/eM6iROBg4DK5TYbr6M7OfDrYzixldwmEk43E69pyJBbB4TovcvMGFu//g
Ul0dqmwZKuJhJVnr3EYuNgJPXT9fVcvr5f8ByU80mjOfilNkMQE1/O5RRZcA
qnrLkA42gsGPi11Em3JP0os/CE9P27jztq6fG8ErIckIpD+bNX825L6Epn5/
Av/JqcOOeASVrVMNGRoobcPn3itpJKRdnnmrF+1G8ihUlIeVlgoZnchWLjzW
4v2Ru1KHLj0gHZovLDgNACDyNRYTXQTuOypQmcEjGR4nW0gZaozH5Ggt0OgH
zkJjmZT+xvUEXA5r5ZPymUMVvJxS9pL4Rr0KvklEftenb9w7HNLL4+hgwyto
A/mOJlwiCOGSHJRhtWJbjUWs/vTvhcEqPqMMEIKLuZka5IbH0LCZ6MYgeJFs
oPV6dHT2WLhPPDBd0jOHJ4zFnQrWQ9TpmCFLMNVXKUwyIGCv/Wjq2cO92Jzw
DW9AyNUsFs41U1JK1GudwCCtVe57MoZVVHLDhIx/yYacASQf8o6MyXLPU5Xg
Z4WSZFTbd0PF/ma/IiJcLWbkGaUbbC8dR/Fo3HnC1NsfKynGc3MiYxvUQnlr
OAuYbQ+N5Big1dPFemyIt1+YpC+qE/MqpqOXHKT0gDSokWGwoxpfsGlLqrZz
bsYflODbeXBI/cfkQ3aUNdd+qaFZit40QMyk/awsejgG2zCNdpXW8ixxQOms
yS6X7xQHh9JWTlOU0dTtCffXHmXZMGp2vl5pzlL6NEJaWWTLR0QcrtDL8FhM
aJ0ZZLo+LD84AsMueAjNoPlidlZvGSMWCi+HBQXIDMOI8qsHpX8mQ5kCrXa6
JKaC6cNXCsobI2nXz9vSIV4Xd9Bb3ZHoRylflcwRt0h6uNpP/xrTuXo4tSdF
EVJlC+toYVwgPRxiVRkJluxxdYJetlNaEcHYZRPlLLIS3urWSyR4bY9frrXH
3eByaus4+zay5ob7FVJ1TCfUaaMMwdoxy59kZloatZ7YLeGhIXprwrVbWOFN
uVKD6beGFEgS4qHmhoYGLP/ymKe7IN5VC0K6wxPO3+S78GPG6bXv1NgyeJti
O+mMSszGLTD8JAtCuVRhyIL4jNvjVHaUBYH5HqvIPyH6SY3oHoX4+hDpB3Vk
08TnTY9XEqaXwwMO7x8COq83uMKU8McaiPiieKgieYnglqPUyyvhzCbZ8ZFA
x7T4t8Qtr+AvvxVkqbe8wc1PoMn2jIjCp0qlVO9lFolXi6irt2y4YrLZifwL
Wflo9FXPFpstg1rJl78H9TNzp/TiisG4tvt6/7lsCxxCXagVGEqoKNjA/pdA
ygswTHQ92y1KTtbwAhJOcdBSbRUV6+9l0f5VOZ78zOU6A+xa2NFp24PNrIX+
IXjVaO/6TEJS5JM+zbAH5QBNcL+8tKN02Lgs1N49rtKrh6MuMCIML3mfhlro
6gQ7ueyUxQ3F+YZoFrHITyELC6SzHaSJbedqeXO6kApPEuEdIF8K/4jTFi+8
wXDMHQMCRdHTAq3kflA2tc4Fi6KfYNE/1fFEtts1cgm0IjJlycvuRvk9mCUe
NQScbcr/PGWV1cAxNql3mH1IJ2qqgxuZxEW0DH75wYNELQlRgr1vsmamAL2m
xKkDV2m5j4zbk8C1gQjX3HCFLgfFtmuAdQ03sAjo6choZGA6yGAdI7a5E5Mh
0xMeRxUuJxYgjdimpsFxCcTTJTivXITseNxsjOH/IraMuD4/E/LOj9j7V6Uu
KXhRgHpZZO0zu8aL2iEgRlhYxs5k8p6+chkXuMmXwFHXZP1NZfj5r+tEBKyc
Yu5EavvMGkkjzcG+j6F/fw3kCVzRvfOUcFDcfu6GBaw9yvigAAgDe2HhleNS
zDCTf4kd/J6bw4nc6on2Xpuhyhcrt3ejZSv4AV5vONqJwf+IhcGhFxv9Me54
UpFRNJY4GIVtgmAMEJWybbEFQ3EFnRp+VLhm3JgPXqijgY7+Bl9T33m8ydg2
SQkSTQzOtPsc4REp7QrHekIw7sXqMLIB+W7BaVSVPDGOxS4t+jM8vtlNo4A/
QTnz84k/cS7XtQ7+g941cEn10IS6mA5P28tWgjvf2hNcu70J3nGBoPmK+RRK
3lp2kpofxm/CnNLAkBwXCIifJEtc/rKvBmvmRD17uqU8QDzXUfE4mr86WCzS
IW1oKjmRXS6dG+sYrfU69hQJtVhgGCBVo/bQrWvBZ8zTM5Dzxat0n/l91/T7
U1s5mt+ZFM4iNOQCBPNakyXPHINROINVFrLGSDJl/kxkON56Y/QBa7gIEEwI
vBC+AoXP6klAbDBTo1YwTQjcLAqx0s6fdsx/dcGgWwqITbo1niwsOduYJDcp
FVqL1hVYw58+gxdU6LIYlbZycjZvu80+sn1bIZFTWYMG+reK4muaykyu3BYu
nbXpKGdfREeWjzjiyCUqLu2LP/eQR6P7iWq8z9yc011URd7KynN2CSDSjgep
NH5KXkH4iYhLvwQp8y6e21bfxeaxvF6uEYDUmE4mE+Dyl367Ui4Vq2wcSiC7
/H7y+G2AdKYnvpGx9OG+Po1fCEVEPW6ol8L5KyVp3N8bJNRgKmuGofUTTi9G
bIcOq3SIk19Z3SaUE+TdhyG2v664eLTjZpnKujEfq89ePf18AJoczY4xUAJs
smnXmEmsFuK2oLKYYZ+jUPAQvQnw8WduB06DEGUUgDHEPISYkfMGFPCFbMyV
eXpyqDkXGXDGkY1JZSA/XHjESfYEh8zVCUl9veUPaz+Jf/7i+x0Te+TmUTIb
1JFJ2ORDxldh+QWmHV4kn6Utt9Xvw9t8bIkuEVHvrKsuz1ZTx6ERSjEsG59A
ZpTmcqES7PpwmY5TOvskHFjbTyUD/DoiwiRbxPD2OuBWIsRIXrCof0aU41h4
h2arOut/1LQTtJEGewOI06LzTDpchCHcYFfqjGBrUIWrMfgfUfYdW54HJ+/a
ft8MH0qN2ShRMD18bFK4XOxuN3YwljFvLC5rWkZ0FTZgRd+nsRhkbVT3aWBH
hpXQ5XPNDebwhT48SRfBSzrUHpn9vGrpv+Dl0P8T2ky6LdARRmN3s0+zRLuL
QF4RAh6jIdBkpzYc1h4YpSckYJE4M8K+bx7yO2fLN0/VWTbnY+B1i5gJlecg
h31wfWxaL3qhGYID4ylFUWhewvPUi4HYSXf7YT/C2cwu0jwZyPFxEBTyPjcQ
hOyPcH3/8ad8Mg7rCjmZoEltR40hXCJk0MFBT6unLNpFzhJ+YchqbOEpNtPs
VhMHuK7hnu5Ew+HxbsdF74hvIN9OeBp/zYSWzokuglTsQZh5TBNIcQqCaqIb
i2nZlb5y5zTRk9WhFpQyXTKDrFzzHMouQ5iZgtSdrnSOkuq+Qabc5jViedZH
uPac39p8QuwUg3WBTYXXAkhTJKQDct+QqkemxmT3oo238nt4qt1rb/MymBPW
EDNM/58OqvLSy5G8o1rzVZ6du09MofAAOS+xDKc/yEebkY2lBYkZ+CGbHJNA
bbjhD//w8wYHSzw6gUxrMgi+GlVQmDrQW86B2mE6y2lMw6DSsHSPktS7NjTC
QmWNxnSkGZ1nDLFQA6B3EqmufiS8XLT0LPaOTSk1KdVJpZy96IQHDfIZP6CD
oKg4g5X+E4b7P/N/GepLcqtJsk+Wbox9r5knbqcEDhckw5v8nKp3mGpRcFQw
dzDPgsw2R6s8uv4pg4B/YUspFBpLSrPogCA+yW9AiSFFqN90RECa/1X0ifC8
VlqExGGzaFh8AzPU4jc2JWfzLqZYl2gQHGqmYsORNXmXTaTUWjLNlnbzLI2D
CxcQWIRMgbOEOfHQBCYoaHqyLh3gK3zPIrAE3aZytyUM2vek25Ngs2Kl5w4q
v+iyNXuhK4MRLg6P197BL4fPYDetmFpfcF1rBnpKamHTnlv5oB/fkbNS63D+
sDi3ypwPTD4Ta59Z7B8Gn3bKBChfOJ/94AMzmp3IAoFEFMkkbl257PJ+vfxw
FaFH3H30m/KZb6TSb0KBMNDLI0MA/7aVNiSlr+UvR9QSnofHuGjZlY2+r7VP
y9UpJ6HB3VjPudwlNkCtCmtg742hK79hzelP1Q2eavbO85Wn8IoWhqssKsXR
t+Qj2Lxcm0lozvkJfVcnI7kNpOagq+D+t+rPLxoZ+0OZgogfPGE5Gb71ixVu
+TZpXGFax/QisHifC84HPKDCC5Q52wohvXnQLnfxoxhO+47GmFEvzKEwNvI6
m2YDwLCsGlwC79dUINA7RRfRjfEJ0R5bvtcXvc31cWHPqbITa9IpbNhqw4r7
6WHnXE1u4+dsHlW0p8wo8cLEKkVzV5vNIEmfuptDf3JWQtT2edqz+CMTJAgU
njcsM/zZoG3nt5DdsnkCk3OkuD7xUjf8lnhKMt6aiCidskkkmmApq1H+xLd6
Ch5WzUM2hlLOpb6AlO7QSddr6ux06qHEWE340gVcvd9D42r1n6yhINNKNoyZ
JTA8a5dI0j4AlZ85/O3/oWGTJoHGatrHCfUsP8B/PFFdCbvWXmn5QbOCrSL4
STv7z9aaLMVflNlZUDpHcnFSQRq7as9q1z6qNMmaTgsdh9zHzeWYJqgGAC+w
JOqcZ2xSsJa3syo+QbyFWtKyIFfv5DIAwt2IZIkHZjAtFMl19lIV54iieHMG
wZx/1fgd05FRHKZ0tHCjmLh6HIXiilCnA9nuKsUzuhb3hxiG/BLg0p3etBPw
soX29hrzmM+YvnqV1GUmfSw0ahgxVxZQq69ZdLS4qVHCnuRnR635QMnE+nI9
zME/ybrT39wEepbuX/fvzx7M6wcn+JH9VtWzYXgdM+46hmMINqC4lZn1mwEe
wjT6x9PWMZPMlCM9hdVWD4/vvwhFG+4NCLvdT51HTlTJzELzlIwLRgJoOpf7
90fjGQ7eX+IcY2sjHLe8Wyb2eUKNzMXL/0MSrWF5Za7mLosXm4MclSV/74eF
ews0cxy4/UX9oubi5ojcfCnVskD4t4Cx0vvMgKBb2z40RfJ2VKy1GOqUnu5+
e3ru0ee2uUPv5/YOGQz85cX6ZVHOjIHh8CvjejBqOckn+hzBiGtJXUUtDhcP
1F1btrBpNtvqAJSg79k/t9EW64bm5nUeKWMNWqTme0Tz3x9awCaQHv45pplT
Jv1oPmBvA98VLWKuYlTqq9OijDDd7yAot61WcOoCjoqtUQTfKV4GTg5TCpcb
Suj/eYQwPv2fzwwVbQPTsp+e3+Ov8Qh/ITPda2f9HKwE8/cJW5p/xkS0uO1o
1pw9f4mmr+Upby1nbNbp6KntP1YJiYVp3JGfySTXTBkljaAcj99oOSRKcNrL
VXPZupWnUgIIO+BApKZ0+qvgWqsiHcrsAXwuzFDCbpHrvkcfN5usbybsKRUk
bLhPiTwKK+OFuIe8wAnGl5GW0n9UTlKOIQzW4L2s1WZI/FLfV+5hTBUH1sQT
fgoiF0VuvybBAMTBZ3Tx2fpeEoup6Hx7vN8mWXdSsKz/cNccf4OAmWaqNpi1
zDEhK0AWLpjYor30GPFd5Bw02Wj0Gd5nCUd65syRAd62UnWrrAnGbOCQxTl6
3L1vlnSderIB7b0SB10gGdM6G8k1VFIeO+M1gAPpuJwhGnW0/Y5wwEprPmgX
Oy9cYW9sh+X/LIn/2mCsJl12UvMzP1voDM90Ue0VkzI+N+AfugPTvnUHEUyV
bToP8O1OZqMPfOu8eGGqbxeWrjPmeNu9vUIgvXWJrHZFTfQ21mrZ73C/SQE2
UwKRn+SCBc0S59lWWLwhvn7X6pkwR2MKl0nw+88plqqxuZVzldRSfsKR73RP
wFSAZPUc5y/b39Gc+wjiBpReQvSzsVsMOSdL423bwnRF5oWEp/8KBFo8eTeF
1X2v61nhTfNkGnLASAvYfGuWPrnjMyvTzb0Qmy2s/o8ypOOeUonVtxXh7SMr
IMvDv+eCe6fdDelIG05UC2AoUqz7PbwxphXEYkafQF1cW0etG572pgrGH+P0
FlsOJdYHuXsS4nHSXXgbMoLxZuf+OJzNM/8LHkZ9IMPsy3gJVwzW7rHuzUyS
mIFvGxpLo87mGXlbijAWR36cCSD551Ke14VRwSoQ7mKjD/YAgld+tPdWeVat
N3R3WdNDvi0bJm/D6ep5RkAjJ2P2Z6DroBUr+Kbz6+cPJIh+ychB+m278xOr
y06MXcfm92CvGPi7fRGPp19XIr6+o/nFVfhyMH2eNleO0c/3ej7LRu9m4oVF
mb/sHuGbr3v8az1Z0IWj1rmM0JnxV7zE0sRFADeyWqPXK6r9ldLfHuQyL/D0
5E+BR8nQbYOmMFLcPdzsTqcxlYJnKQmUgoZTClcngxFlwGOQ36i9/4sBhR4U
T6gye4UinzvjD/phlh8YHZK+I2GDda446zJ5JWKw8rX4O6j+0YkkBqeia1tI
v/i7zUhtC1wjbbv1NP4mZDANbGxWLzd5vbMKLDHUiQdnq4+QtfzDRvNmndox
OcUfCdVysL4DlaXmPq+M8uIiR/oj0dqslV/gkFe7imsCz3h6rQq9Me9RorDm
miVSDDNZy1hTl6sAQcI37hccaCL5RqwJzpYjcf58sjO49tGl1SgzTrzZIzOz
nM4kC1x8gkOKimVmRG8+gvDKTz54oLKB8ZsFZ1w52rxgBr9Ugk6ISVGtScmQ
Qj/r0Pa4GXdJrM91xHy9Tkb+2w4sjd/DfarF0U18fGdRLNDtljXMW99zjm5p
f7hoD+i0gypr972VHtyfzMnG8izQUNJxmnz216FvojS0C8DyWIFkSD1QkMT1
e0xWTqGVxJ56Lt1G+MW13DeLWvig2i77pBSwgShsK1T+pge2+SkKVqOKBpvp
x4EZYadx6kBRXo0Swk3J1bAv0l5nMgIqq9sT88fePCabZmcorH+73auiSVAB
rgUWSr2Zc+XP4xIS9jl3iVh51p1r1p0hPQFFqI276wnXXbXBFYvY/tkakqgo
KVmuy7FZqNdAJsiFbyJ1Lty6C8on0PnNakd8mU+6JZtXVcFfAQ9fFmL92rLK
fy9WiXsitJ5M4u2Q+F2y6b5wMhry4AsuXvO6667tCgz4VE7ag9qaKzXPCLcC
JTHPCHwMWTf4M8X85u5E471g7N/qeWURFG0LgZz/j9WybBAto+ZHNa2iIRSK
a8pzijmVTvaejKe10+a+xwdRwlLyrsuB9A8FjPGOKWOrJL27gvfmH6ifWh8z
od7EjZqaqEkU/GDQfq8jVGaCX5xsFlbuzjsq1cVjcYHKowwVq4xONSwhIXxv
mw50p15T+WRvrzI7lKHjrwDbhwGKiprnt207z813E2tUvH4gPRYW0nfayFVB
IIafbSNzacBDEU4F2uHB2zJyTvjAj/SKjlCYyzS0Zu7szCdWSeJsqRpIe+ma
J42i+2AZkJk8vdcysOv9IlE/FubnerGPG8Y911h73OwcixTwgpH4HYXLkbJ3
uy0ArD+x1/B2WPT1OMxKMo9H8eXkDn4hmqCiFRRRviNEw1207m5yebJuY6mT
h6wOhx+1ZJcCj+zT+gI4k/2AuHajK0z8eJ96sXebMjYnY7Dlszls/zNkeQ2V
QmDvqumzvB59pd7S9cHgP9Hrce8jEAYmFxuBUFxHsY8tDiGGX1d48Swd/8tx
UeNfFG5fpICJnCDQfwAlyh2ONOLL7ZlJuF7uJM/ZlI/BEbwus9jGy9fN52XU
pEIux5LuqrapzWfEmmjfc+rzxl5OF56oIBmkrr5GhnQIqq/GGhrM/CIxjNHk
wKF+JtJ09C4tZpi6+m4Tisrm4ObhY7jJUTSsUvf4yiXBVIehYK05E7Dbt3/2
5O+kfziA3PCuZ3l3p9k6hPyYWJOI0eM8CDMcBSahk3mZIBF9TllFYWG7YQfn
QlyNPabiSBTUihkZLT+WybYmjY2mhiUgthT3Xi7vWrauSbbGz3jD2OftgIcE
YaaKzv7trOx8BYVqf0M4M94XO6mTuKIa/ntacw1cnbcAfPMFt8tUA39bHpYF
QJ8zPOliBT6O3LgTyPRkoyxJj2N3UByozFJUamePNa77ibGC5nK5n8Q+yJYG
jLiZ2+IDJdpsZyeJvRzNlrl4K0AmxNLhaDA5Gy3UdoSiS4XZ3wUoIRDRu4lc
qV3i9zR31UsBoHJYUXkGw4Gkh5EOSiLBOvF89O8dU9IhLkaF9yTYm81fTKUJ
FLp/0sdFSd1z5lPfSZAsiYOehp5kNZ9oD3At21ht+Zr+dPQ9dUJcKzfVW2R5
0ub48d3Grj1Nb+T2M+Y4EKRpGuXrrBXCqpXPT1D8b+l5xz1R+HkNWxCPF2C6
tTVlZhjDFN4ZjMycxBmfBLkfo0Bp5jhN55BOXD0Hl+0EkR1ZQedXP+rDPtOU
GBIviEIVdCIA5MWwsDYOEA/PCkVpEu68cLzQBAAuPzXE8wE1D3ZeMdhO1kcT
gzLRbln07F1qHFdptlJS3/WriNNbTWzW+UXVTZQcM69OHalt59NK7isgwtku
2pcF9pn44qnxv48rs3k/6fgOcjzxuGRFrAgoGzSk6tapbh9ghiJ/IZcmCx0T
UbBMQ6lBBDoRAqyD7tHSZ4M53sq41eBjm4JLv/DF5Z2K5RttMftf+ZkIc7kM
7z3E88aowL2cnGS+wgZSKQff2iEaVQt67to15019wejUvwaw3w90963bUTyb
W4VBPiTipHPts4VNJR+kzsZG6fuQmCn1jAYDp6ggBMO6GeUwpslFbaAhmA2D
mZPt3fT/wPSXr83UCNU/aELqAE+2vUso6rWRap9KO+t8f7Lm0vpM133eWpL5
SpmNZiZfAUltqccJ1rIjyoa6BSwH3wHjoqkLN3MVxBmN1IA8ABq8gnpbFnxx
gdAcHCztaRqQ/i/8dVylxuoJXWXZZKIdI2mIt+PLJhPUmNTzMAxea/71zNFD
M1XJwMYcywLlp/cffyKL1u7b1+5jcBzwwKBKer1RTj54gkRsrqwoECYK3ann
aPw1JLneGpxwUjptVrtMENmrzB7A6Tw0qulFwL3vydQ1QotUIFWi4AAfkPgu
3kjFaD2b9G+gtAJMet69Nu/piNDaFWUqhRbUc9GscQVCn/lZXvHFMXArm6n3
aD/rn0O5S832LEGfgwiB4ubPEjG1DluYxfcmAUpjqxV+Fxlknzm4sI2mxdCn
By3y4XdUlOQHLnQEg4wOtVJL/STJlIRdevpz5mSqMQ4yzPiL+FbhiX6V9PFg
GGzoNC9aqa19aqIHBExwWJfvRRmluvUYlxqCVbqvKzfCUqdcVmfImVoKRvjy
fBAFCwBGZO2x3gdz8iPZWXBGijXRhRGcpHKbRTG6Z7t8bYgBjzpiuIkOsKCr
yroUeInhr+eZP0/Qaw8CBJVkPEnE+ZL5xsf4F88zChpgyC/HpI0DECgkF75c
ZfOQK2l/RnS55bFRjt5oRbnmZdSWPCiTuz2Z6lRbV1vCIZ862+vXSEGeZpBn
Nd6RjEQtaCY3reilDPosEZxVObzD82yRbl8F0o10cKC+zhzORUsxItsZrON3
52oG9OuyX4BkDUgWyL5pTrbCj71LtQjAY0l46fVlGZGm7oZYV3bScTfZAjw3
SBmYDGUBLKvZDf1j3Q2ja9XX3ImrZRNC7yXedmF/Z5Vgt0vZKN7U6dzJxv7+
TogjpUCuUD84zS3MbXm+mFiYjVBEJeNrdRPKuwh7eV4xuaoqTgN4bhlfdLiI
P4H3jI/n3+Pii+b6JnO/naFollyh5ub6JlyBFK3qis2Ra++t7gh7aDZuRz+W
zXS2ovO7LINA8rn2HesIdkatm9xefPlmzuYIZifTIkdfQtxPDC27I8sPEwI/
OIwCvouys7GOSRSN/LZ75bZKX5l0LoQ/n9fZe4R6OUOLVDYUpK7D2CKqmoh6
aqQn2Z7mmHvdCdYtC1+NflMp5rLwbz4gaDJMldLymGT+Ajm8+nK92K0Mu/9T
O62GcYL+WSP6hWl4eNxSfMhPUAZ7VlEs7PCgs6ngw2D6Cw5P6ghSkJygbYJp
OVqVyW9LQRKe+y9zrIGVlnP6XT72HL09q3fytO/KtzXPW8VJGCKPTRFSOlhK
GCDCAhUGSYTuIrD/BV3IRAuW21hTOK2NE1gdH78a2EdCD5o4krunHCUClhwi
5Z1b4v1/VeLEJKDInOnU9N+TMcvSg1V6t2nfssKH8YEhMzNs/Gf+NqE2YmJB
qDfYc9KMqYNLs0uRuVNLhjm5JOMkn+TbIUf/H4fxppBMhd6+HRkWfCJQuKJG
LOl8nIpTf6KbtlPXGDTO4v6GdRH7BU8gCk11qXtNhqC4oCYo3Z+r5K/Bk8fX
MWrP/veZJgjF/vrjMOu4zTTzz2qhs5nW8jgWErmlqaJkInvkO8baCpkG3Q7W
aHi92FRXFj2TiPbFGwnJHFUooMbDMJPsKZzordvU9OGWGYoreEAFY67HQnkY
lFujrVnWtKB3zQPHVhfu4w9tWiKASWPn0wA0K9pg3p071O8DS5ar8rFyn6dq
sVhRvyvSzvZdNG9qYT876WoMIR6hCI0AFwUZ5+a2Xhb+QlBcVwVkHZbFy5cE
9jvjUrxAiVQ6mSk6NkLrnZBeDR8zMPMd+8g7eA0EH/pkpJNhjSs9N2WqSxbT
IiqJQ7/K/nbybDqaV418NRGjMkXjSSIxbtHGH54i88B8oFu+fnHsdoVHckTg
7Fhag7Um33fDNRzpad+1I4dsoTpFo0+G4uWLvtgGlFEjEV/UUsPAo3Ym/n5X
NG8mzAFaOvLLnkOEUgNn4s5BG2iHVeC5GSw4O0C0eZFSwucHkDAncp0x3NA2
5VQtfMrDshXXcXuUfWQv8lDJLCDfKjPUZFlBBlQTIU+D6tYPQgZiV5CuZqck
MsHU7fIoYDHXMoVbJ1vji0jBHwbu2HtzveSnJtrF+MRcap+gzQNvpVztnJKd
XGx375Q7XdO4tYQJM3raw6bA70+Fu+Wam2+Acili//4eZ+2IXUU4G4281YQO
bZGXg4hVzMP1r+2A7Ba+fUbv0hog9hO20aMbftZ1ctZvUaAm53wIkVc53BrP
AoUJfdKL+RQQh7PlhFZZZ9wpo8hkPp6MjyImDjhtl1gbwT4Ihm80v9hGblGj
BrKujctQa8F/yirlJ3hGMagr7moExSwkDDR82ZZ+gMh251mxPczEZRvNAa1l
8TzBjRXguRUyoIHgKD7kLdi9rTUH5xyhOTxFe7r3navJIy3a60QhBQwr5Bcr
05007Tan9NWQyLTral/mvi+/969EC+UQwSUAKUnptN57rqkWBqLTusR5WWvf
WG+F5JvcNJaVMZ5GJkRRnLcAAkuRUdVMpPDyxbH9BjjiagZgYQdEdmqXIGOK
hAQbjje4tsKCT3Ldf1HocUSWBZSxcCdRjbmg3hwVYgCVKokiKGTfpCgGmVhL
+5q3eiuKqNo+tROAIOb3M51Gbhc/+XnBKMMfI30WlKt1ferWbwtTF3YN0WxX
K7qyCrdsxVJ8/D8VF2ieQvB8w7a1amg1LPHBDGgGilMD/nCIoeXbFHTJwdgT
RpFX9htZcDQnd1YOlLJeRDUhLdxDj0uTcDhguyPFOeYNXWM/+/4V/UPzxL4T
SBG+FPt5SgWnWdmYdzGE5YwwgPpQ4E5eb4SkG0fhC6w7UX3zglh37tC+oUHT
AMJ6q4ze1yW0z6Lf+uYktrxM48DpjzIO8xb4bXxJEcwrDq7aY6uJ7vSGoj0q
paSxksp7XW91pMnhWVa6/s4uoL/a8NlfjvBW/M6uua7qfJhHcWB/xjIAZHNs
XJkqnKCsdurU5teQ15cp1ExOADBw+BOtM+fG3z9cpOIevNm4GgFVucw45ne/
NIX5WjMJ8P/zESc5AVOAkZsB0qzvtM6xnAPlRX5pZganqZT8BJQeQOO8asR6
5BrLvFOt9fWUK9+Pc8M7PLJ3ph7vIg2PWdthpf3BNpyFvfYOjx2U4GIywU1f
sl4v5UuIFvi8hirlnJdBAVPE/qewxF7fSrsSApDeYUfmotA9Q3RpLd9ArEsC
YRwKGdKYqqN2aMvyHFELmTE+NpridScnkkzfdUS5plhHpVvG9eNckBM/lGyF
PrJkJWjT/D+P+5YghnbHgiyQhxVHLSP6LyTGN+JFENSME8f2oUDjp+2x5MdN
W/x8rF40vTqoiKFAAKybmZgEY6dt8kps3aOxRcSZH2jzB9f3AkhzyfhPp97T
UhRnQtmA/lUlpyJ0qObVWs2BREW88Ge1OArJQzyTagxgagFlrTlYQsEqxHCU
jw1ALHFZ7guDVrfIHuLNhFNAhavG0kwkyKw8UNXJbhjjEu6f9cjos5WP0EbO
jEAgA9sft9eZ5UaZRbpfTjBiWZ2PJExIQvz4cZMB0Tc2EPKMhYeXtK7Q0Y3s
uG9tvR7xL+Po+Q7w3nAZLPdrW2ydmlm84SlySFq/WbAPcANQx5Ej/1jdhP1j
mMMMfQgXmA8Fen7fTXS3GIxKe1GH61woPvRli29QNcv+QTQjE3FvL14SZT3D
vXPftJTWk9xWGZi0uhHsz5MtY8075lNr34JqiVqaJ1cR5tYaB2DFxMtNngd+
bnkvP6x7fNwy1bsqoLuzdpxi2N6yqk1jhfLI1UgGgi/5b01leA16HFHwAv4u
UMwZEysdB+T7lNA36jYyWV17REFWFqEUS6dIhSvYxJENG93BgCzpDmj2nLye
De0EtrxCSmNCmQbN8sK7jUw/XZ7eXsuQPYhANT/Ycdbq4Z7PDF10xaVLUYz1
Tor0Rm5jIutQ+C+5z0B/qxcUYZbti1PK0ZNSQKWCRyCqzRkpWM8dG/cABUSj
OvnTHBh4UhIyURMxNVSCXTIrvgRGEvffMDenlsrfL7QaKSMaJ67xd6OYl9UD
K36GwlFge5ZUV+wsUYUPQL4+epR5C5b56mt/RgLMG39fXvB6YcVyQ5zHUq1T
MKyfQ2uGL9/8DZP4Jwpp0S2JrZs083nR5tnm9gVdFKrjnJXqI8OEYIv5SNgA
lqJrSHCrdpXnHy9xptMJQX5vRlzmbsLLcRX7lWzGD9nlaBI8Ddaf+kz/PXtz
XQtZqwZa9wqL73Jq7RQLkyxH4f3bajnB01Tb1pc0RRAcYWyaX3depKod/Q0+
6U1GiJmHXm3WiASCGMAuP+ksNfEdbDf8k4tpGMW4N0y3uQq3ft1YbQkXRe3i
Pp2uxWqA1+If+TOLLOuz340Oof0KuRdcPf6DvDOsT0+MhCuuj/SF+fpFQyUv
kOVZpsUaffXrVbl8sq6lt0pN1Y4zhbt70BTQsda1rW6AZRYCwJn6tadzoE3L
amiL10VPD8xK0qU4BcSN1dli0MDutKEbVOC3sayIH8PTpFD/kWFjv4jA3pB6
1dFgvVI/nI7Y9PArp4qGadgKyiu/ky3Ef88u3+qXlS1x9cX2HF8lqNfi9/2H
kUjELYc70cyD5TKsMJOllvCWWx2eiVXripmkj76Qf+FNr9m7DaM93HAfvnS2
MLgEJoPZiXi5UDEbHXspqnofmo2LqorE0fmDOjGYTXdZPstNkYatfW13x/ac
yr5rYMYGhvpHG7/oWBj/o6HpiPYGITtMkwNxDc4ruo4kEEAEFg85Pjp3c1sm
5VbyP0AcPRzV6kstQ3xhv/QYb1ZwEf4yCAdLanhArJT117+eiQQNHWDA4onp
C9nim+6h1GbzY8cpt2T08CjkCY8tSD8Us7MDRe245NQAjsusVlhsVcpg8Yat
FhrVSVnftRLPwkC7V76Rd2CS8YZq+cyHSH39m2ZUpdlcBD5PuBH2VgGVqfNO
Mo9RUqVb8jaCKe0rlgMgaH95T/OiOompGqXQbq+hiInEni4a2qKPnyB2z/Zn
2SC/iIL5grNirKeXmaOdPxXSPvyUVSCI9g0XlVHv7I9Jf8CDQqloPB+mrRvH
jV56GIOYraTb9v58JXPUOzGrYbfhUS6Nmk8L7NYqclHylfQnWF/DnPV8s7lv
LJpipb2P+vkaN3vC5jaos3bfzEFNQ8d1zFm2P76LyaWEPahHX+ztReJ+sr/7
VZvOBuZWgygJtzzhWrcCfPFcd/UN8ryDe+GIyR1+wwFIe+eKLyJro/AzaKGA
Dj2lbUxpCS4gGUN3h3yA8QKPI3TVt3JYc3IpfYqjJjiN8vqYJ0nD6UIJNXxy
6/cdxVA7NLN3T/t2iPYQX5nC+11PeP/Jz6POfnYqeCSAdqJnEpvt5zDB5g7K
D75uNJ+F2e0VwadyplvBPVI05+RPF1pMAjemENVizMDqS96Cqb7K2pDxNLfD
0uvZ2+sfjlvhwOb61AzDNhPfLT4o2jOss4RdjD6v/hzrSxsncuaFoRTbpQUA
eKETHahveX6qzUnRmAQ1mzlthva2aB0OPbz8lF9OAULCYKaDqMMTEGS4BTML
RqeRKnqbXeSsqjkatGpQr/8+HdVWI4akwhAi765qD7awD7Gwxrtkau8dT5QR
tvCjBi8AWZd7PCi+uRYlbaZOPlL0xZrJlg5Xd0EsrOiFUqawKk6mGHhxKMDM
i6ZZC4un9oQqzSLMTRAttJ4QsVvpL8NrHDOlQncIqOh2pByTWraUCUTuWiOY
1G9CiSWyEbbOBsPrkhoV7BjBOFpSI61k/gGXA5IHPsRk7DmQVV+yfVg5y0E6
8KZA1Iqztr6LIYmgz7pSwl2TSA2rTwrT3U3rL4tjilMY8cuUl673I9fGqJNh
00fArBE+hsmE78qcp0S9cBE7MN2mtIl5Il8x7MbaSLNc+Zwxlq92+/mqPVJC
qY58jhKNDPagF6rGX0E4NQXG3CLNz4ksFgW8/BXnMXFLO7l17mYmsSzaHO87
X688LZe86ExsNKS2CMq//yf9ooEOKAc222V05wa7uArefJ4hqM3ocYfOnEMD
WE2wjEKjHoGgK8SKQEabgRqUih4aMX9FEKw1rOQ2BqSECNo30BiVigynERSM
VKa99M8SD1ViiObP/fKJu9I/KtD1Eh42SGtv6/9P5lo3gygTcnGz3v3+ZveX
ayEI51ZgSNqsGYksMCTXvCTzUxcGL/kGeOuErO6cVixNnwbHNqs+YFe0f+Zd
nLr4e1x+DnegfV5ivewgl3dCRNTDPpfWu0d+he3or9WPJfMtDPHFbrIH+9GA
F8Uaa1SkrBlcXuBt8p3vytWP58MQJwsv3E8fIA4d/j4BRii3sEV/EVahLRCc
RPGiZld1L8ltPrrY6IB/PSRJJtVKSIwq7em6Vi0O8+rqSlgVr7Uxl3ABVwLK
uCaBuSgpi4L3pVJkNMrdhY4v7ZD/EaLRIErQLudIE+Be0QpkI723+yzwwRPw
zWGM8P4mYMEYdySXrQsCOcvmhcRrKHzBjQNiZEQO1X9iuxAmLiZlLafThnWj
6rJ3vqBaYtKKAh59jjFCqAekSCE8psmUvs/jTOIPmgicy7/asFjodJfvVClN
V1tSQbEofg3jIPHu4MlxZgzMSGAl2N31JcYwNP7m/MYGhj52DNybkE54TH8m
xG4XxXeXHEG+iwSkgaNUuqn4t4iY1rhP+E1dJYS4oF4yer/17G4mAF6pvhWT
kGm9dPX2U4HPokQ9/B1lzg8UADlerVQyEHlcv0EBwSbcnzVvfth4kdjiUEZd
GlZvcAwo1S0rn3SVt0e/QBNT85AvTa5ky/Hqhq2UOhhQn9X+o0U6bzI1yTD8
o4AbY5gAX7lk2P8O06sZWoP7Mi6cbAPySplkZqXKrBm8r9525E92uOotyukx
6GRGUuI1vb8yeFUnEvdTreNH4zRoCTwmp7dHLqVlEvIXJRsxWcMFTSRd54NO
BystyN8FisV+z/6Qci78VoG/1agG1xZ64psa0+fg1gWuXmbg3IJDNZ8jL+ub
4woUu9kCqEZDe+ve7Xj++ZC9f+K6RSyCGNu8WyByPnp9JfGj3f8jczUxB5z1
XvWcECPBlCfLPyMsuw3EBLUnGXSAGTzCJtSqEMBCyRnj5l9WdlqH9MF+dqqa
fibFvVy+jdmtfGtM5VBfuZ67ny2vlmaYG63Fg+E7e5wn6+URk96RgHwce7CB
9tr/ntQX/SvYp3+9exxplRddOR0CaPf8mo8eCi+eMWuwCrP6KmAicFd8JGYX
FRUJXc1fZT4DM8YmfZBcGLxlEHxPreEWloE44QDBlFZhNNUikbvtRcdFLi1w
HQBBt5NII+mlu6mHeyEOAWP5f82ZbADKrx05V5WaxuUE2nuJcv+bLHBHol4R
x6V2a3n+2V4QU3H9ZqGojCD6sv4ATdqYr33mmPAVEfWsuH9zxnv6pNAbA62A
uo1o8Su7OPIosgoVMbIiCsSip20U79rBNwQgX5j0U3udZq1f1D+3lodCNekn
5YxAQISyP6tS7rDvA5wR0HgThpj1gfs5Gb5Wrbs9puIPm43AvrfU+0von2Db
PZz/pxnRrqSBQdVZa3xTpmxfPP8TudpUJ0hhRiNlFACMB5tdFksIl+d3FCMH
LpJKz4vgpxLyBkgpezYxt5JKY1auZy7uM5O6RZZw9WsxWYxo1XnlGLfqCEKZ
PpdxC86psYhOmTCJyJt8M9KsXzEJITPLEBSL2E2xZ4R1q4OIPEvDqHKDqPGI
bcyomDPMkpexcNu0KeP3JHrxWoRyxBh66il17EDpBnxMqrqeCwyHpJ5gBK4C
13BI2+OPrAcgfh+WXi/h4nowUZdR5qANKNlTZXIwKghhrLNeCOFdgr6AtHvC
NRkUr6yn9z07TqMY9NGaGjgLJHmi/WDA4g/PKHZW3y58l20q/n2xpAiP0hvr
f4iML9exzco+7/WGaa9W9WDzMJv3EeWkeJq09zQnfT5FaEYb7VsghWSj1Qxt
T7VhnogBfoVNp4iKOAT4qUBFhsRIzBPaN9x63edYmZqobzTfhaiDeqQ7CBiP
mp80gHGxgSeD3NO+Ai5IpG+eWuLuB9duTQbZKN6Ck59NgptARuWjqwwAan/B
UCvkWKv6Y+S9UxdqR6mKKSFZllhI/n5a/Q1ofQVRTPnk0ER2kOKZrl8CWjJR
+Fm9hjrYqh5mbyT1TaTjkdYNoz1pVMCdOsaMWzBp2wtoIhzajvrq8NmrL20W
BjSvAVZ5dN/UcwyFzYFv2URK8O5JFnrlMbmFxc7gBYYKO1XYvuqxts4yvOxE
wpairwC7C5r+z5sDDMLBMd1IarBmaiszZGrWlFzRFlrJiEnFPabIdSEkLdpg
FsQ9tDCgKuLvYBjkrAb2NxDiN0EFZS6CY2kR4/NqFBmk32KNxrFzqZ9kHPys
bCKfdcbl/K8sw1LfzDHvEiZ46MVBPQAB8a3tbwGuVL75fy+e8HUOJ6CbgTIZ
aWqnjpVD7nYFL1d5Tz/aOfA1QZcSOsPKHWEYw6ha0EnH2NCqfIsRmWkUssvd
xWegiUpbyQw0rCVOKSi9piYPsy1tKOM2+ALBpLNaIk7ftwXFnliPpYDsEpcB
UsPIQKwdJmXXUUlsxqAeUSB7LZQVR1duKvD+wUWHsEQjMlOxKj2PMLPk0v70
wYBOSwXwrdGmtrhE55KUFryAWE0RihDHVMHHmjYLk9182c3Gg6xvUT+H8XVr
fHaokFmyZG1w2OZZADifBktMJy3qYUjfFNgNh6R0eGgGDrM+gUVHq5Z0ny2m
Kgz3aMjVHMRtN6q8HDWz2eYWvTF/TC/+oi1+EzyhEEwru6Y32RvVgVqGeV4E
1FUi0KiPt6JZ8IUb1GKIXkknxiFHLd6dC5yIfK+Sc/cpRHivxYEhMzysZwOj
OoPlMSbn2BJfV1PB+CMG75Mx/wmBxrcGyP1+FkjHp4hj+cHTQLBIPC0KyBlF
9Ez1wvjlyIv9b+Lc13UOi6IwgJ/lGrCMVraKeUzK82j/APkNd9S2323k7mYf
nQuXtf4r46zmneBVfxXqJ346snJ/ixQsVP8AS9Y3jE2AVHam4iTD35JeJaTw
dMufd028yJZVYq35q3Wm4aBarm4UsvfivecCs9mrTB5I2fNxzuGjInAA611f
qMwfMb75m/gOhujhBE4wAUCMBlIi2+MuC7MU+nXWna16XoE4AKywezlFBlZ7
Olhdg9dPNKVfbQu+q90TKFQWUw6nUXs2SFZAQ0prNewzXyTs+gy1vseOHWu+
L79sC1gwCSbrMkZvo5AQuVhPjfKRBd9aXz19+56PEf9X/NhuBuYm0RUR2cUA
ZXrXiV7/5UlSTk1iPkS1eZWZ9vxWQ6khQbiE+ruUQv0x/vtqKHHHxoDhvlDP
B4nuVzV1R2w9AK+6I6m2/Ry2eHpxGTSw3NkbfqS59BpTqnvFdwdcei941Zy+
kKh7Tv93m/WecmNCv33TJrx6QRKa0IreyMkMBKLs/+8rv7a7soEtPLDrBLbd
gheYR1PmnuMz34IfpQsnPnPyFUVgzlBgiPu50u7eW0/2PJbvOvOB8bePCeHX
pNeAwM/MTbDuQNUg68qwmRyGaPObHQhQJP+ZfaH67KzLCuj3oZQCZRGphJhY
65ZM3TBCjgE4Qh+GDKoRmjgOXkqjiTthUR2rbZr43PQH1YdC595L+34NXpsn
xyHv1FFyriV+rLGo4Y6uVUSKqgnE/KTepHPHlGXglIZ+g8F6rjwUtEYNL50V
mtxSUmbAZdBdszpMlBJuVPBwlQdd/8SJ6wL1Jre1P0fu+Fw/2tG9kQNzq3ce
lVvYUu3JsCrv8NiTRetsnaCF0BSarBvebjd68pxuwxy2PyYl5Wvf3b34POd7
Hb9CRNfvq+C/6yipaPv82tNSCGhpX8dsui/omayEm2bnodp6PzAu3jTRy5/o
TDQaCAmRDEjVd20jAxVaHplAazB+BPV0Z0OODGBMFEiLZ78vsFSDUtiJTwef
631iF8s6tMB/xXyf8PMKDJoXgLjhyMRJOoIRgFl+46aK8HjGXk4pd2BNcTez
X5P00jnE7F9o1Hu8t12fB0loTNtzuCZPpvKLNMeKITYXQUEo0SLWM2u6pvAq
lxYVMkOCt501PRl/bg0YDQKj25m/HCTShnTyiu7D+uPQHFe8Z2hJGiOUaIJh
jEL0MdUl5G3xfdIcyqH2R6PShET/g22WBuISUWcMw+SrBkH9NMCnNcxcwNtG
B7x1tHR/XyhQDVQ01eygDcNofl9vAOYHzMhUD/Gz5CYflM1671TEgnFb3K1j
7x9j8ZIimXPXY9ULkvr3+zQ4tAEvPohtgmIt5uo+xTirnMCf+0nFkv3MAQAQ
YYkKyEtef1jqDUGHfdEedP3i0Yn0nrdC1t05+SrZtfk8WV/iBjadlBwHpfOJ
9+gWTnj3e/CsZqUZ5uCEKXgCCPjXbO81QB5o7BwJLCnipSkOZ2gVP5nVjhav
eIVVX0LrIB8bTH7O1b6sWTqLA4/Us/R8ltPcVPAdchchJ3jS2NzVCgPn54Ei
ZWCgcXu5Pf1pY1DFvAAToUL6s5kgBV/InhYuf3ehbccKn5TwuIWbg/BAiIvr
KPNzOf5UlYjJq8Arug7VC2ZvsZYhI2hTvU7GGWlHLi5r144SkBYUUjW3OZvA
S2+LZ6skVhd3gTYv5IQaGg1x4NrO9+WzKNg/c5HUHRyQEHmGZjrcOeUu1rKM
JSLlS0XsDjdUxMks0y6vJq8i0t9PvUTjE4VzhbIbkPbChPOGtUCcfO68FgjJ
CFTlFTJXRJ2LKz7I8wbKRJ6GhphjmnM4hv1vIOsyyTXnmfSo5UD/ThZU8M7Q
aYAmVBzUbMapNA3WzCIC1JtbJZSyuZu6Xw2MzISGWeNo9zy+eiRco7vJAUil
7U37WO5WHtInc+kwS4QyjNTOPhRl6HlLVFC5c9M5Ly/qsNhGTMPsrd0U9wXE
fRmxl+3oSfULrcFpKb8Gl7PlxcSbxbobLil74WtK7kFShF4EzopmQaY5dXVe
zxWbjo21Cl5f3VNuUTQODU1OEk/ot/Uf2jGVWN8HiXy8lUfYmYT4N+DBWor/
Blb7AIjt8TjS0UeX6myKIJP6lna7tN3g80PpYdwenOySLOpSROVl0N949n69
16bXxQ4qmaKg9X889UKz7tpHlseXTfqdtLONSOt3vT6Is60F/5c/urE7vx6R
xsS6MQkg5w1Xd0IM5yzNLNqegePoQd0NBwp70iOQo1k637Vyu1hjzvgexDnq
3zFWHS/AToxgkq+6slUw0iHGUbytLbTrQSGjVQQkIbU5jzF+ssvlJHuHPRKg
BoNjQI4VmRk4+LUobxP91YZMUBjjxi7Ma4iXzzT6RjzSr5vM2IsEM2iF0b3V
hUtnQ6OteuIyscBF1HmRF9+hL1VbYzZvA/qpmqEnQ6Q5s4bLe7M0bFMqassd
JRUZvvSpJGffYqRir3F/JmKAlMck8F2ld6GBdtJokd/kYxZSf3td7tjoXE8Y
ToDaB+ZdY6kbR9WS/ZYcWuGx/GrP8a5NrYw5vso9MSF4yt/og7SBG5YXoflJ
oQOrMCa1MAUhB43IpT9M6jTPKYAEad/6yTUYWDc+IwN9zytlrd2mFIaLiRkU
KGCeNHj+RphvhQhIxCWReU5sD8kyAgIUaSQ2yDnfZaqWuJntfM5c046f2eda
kOAo47NJbuP42PKHlVAoyQaZPRBjyFCEKvWIrCsB0eUvTXwqnZ7P+xCcGkZV
EgOkH4cuMtV7aSPi4vxOYiosHXgmAXvMd3tfy4LvBQaM3pYYfuR4juHQnxkC
dKai/4AZuhceRUi0saQpK4Sh+kRK4l40vWRvI/2+v4P7CqdbbTVcfgvL+jAp
mvRyEFcLZiloyvJSOt63PX7q2elhWSNO2TyRm2wIzakm4S9PXoR/5/yNbLxT
H+zL978d15//7dVs5DHB4oUqYTBTv8D9ffq+VspAyXRY/0/6ZypDzPo/W6nf
nRTWnIMpxUf3BUenHjiadKmZOmn1CrC5a4jJOyu4kMrHg8cYU1CAbnPGM9zG
xStTSn8fY4PTcD1GJRlJQtTEynOyrAMmYueJOPg1Cw0t9pdWnoNX2aRUwKnv
xxOPL2M5lkNc3wJ8Sf4MPu1Myi9oqn3sVC2WjLKjgZyJjKTtGsLyFjPdQT/H
lz6SHmAso8EAdz+EYi3IXiyWdgSMRByoSvzTKYX55UM/Zb+INIkTY3KWLB4y
PMw2ZnZBKwrNJNgfCEvdwdEKPHXpyiqT4riqwuxgnn3MuSpVznN998K6iI80
jhrpVbuTb6wPcckCzn8NDQ2pddw9vuSrGYge7qQ6xuGZ9onRYbEXP1sztysa
eO6Yd9ol5o5LK7Pg9FL8WnDmjODhaARgTYgUV2QK7gUova/JkZVVK9xkdt0E
tfFpqO53N+MfHxfnQj7go2qK5ZV66TFyf9a5mkv8FKJwFPsQ/8hTrSUu0da3
6j3yBiqqYU/aKNqNTSNTrix0ULmh3wA+cL3/zycpK79kJlSZlhpVE3AVftmA
U/7mjvfWjBgQ81Lyt3GaS8k7bjgzqWs3MTUo9dukyzC81i6Gcn7EXoOqKKdy
wMHz27kCdgo/hjNj0QNUeha7wU+MWla02qI8Yp242wYmmFyPUZhi6vk41RxV
D+oIRDsKIfim7h69Z5/EQhTgdyyW+e3g/UdSS/jfu9wVC2O81TPjI/H9YTJB
iCgwz/pm9kjxJT6GpbSnFvrcQxaQURUjD61OVH9D8lM3dtM6bFrPlU+8YVU3
df1kh2OFVgcrlLTcy6yLUYP2dwvJYuoZ6Hs/o4bVzn9uc/W7mHeEFB6xTqrN
a87UIdnyei5h5JSTD48CbdVeILEcrZd15LHamCaZsDHpqWnE81xLkjQAfPVV
sy3crYiwz9dDdijCSxNLrjD/VefMjkO2Wj888MsIYtT0egLS5nWQUTliuGKJ
d5ZMLGUMp6Y7P7e7YMB01TRVFK7xz+ORT0n5oecdKiSNxAywR/cGdamooKfX
u6V9DrBT2KNr/TOXgb6ltvY5l0/Zy4nn5dJULbdaJiw7myD9XCk0r9S3hkpb
Q94EYz8u3G6u1pF9v1RaWGkhJAHmw92Qdjtba6uJQBtOmzWj9CO1B0CHySI3
ia0QWo4df7bkkO9we5qhCje+VdQzjK2loGipv4qX1aqDobjwiAy4XT/x+UKj
TwPyXzKEaK/m6f2oTbLWIhiD7RlE/0zcq4dc+Xy9CbPbJL6O4OrRYLdZsaqo
o+6UAdg5FpP1Ps1uOSgUF1/zNjFeAP+/A4dPDe1sK5CAdH/UgJGqGiM0CUvM
GesNhV+49AmMTAl7rJgsrMulKkNTiZG4uxBmmwnTts1g5vwabrR82RkTpPIO
JQqVtphVBebGvsP/a2dlGi+c/6OEPzz6ECEyQQD34VML45bcw5zlhc1GK5wk
HPD5G4oA9v2EcGE62y0v1/wvK7Br4iPsQnu2+paRMtTcn2tlqsarXj8+rCU7
hr8HvJHOqT/6bsTVySEBjtitudR/S4tgIsMW7ryBWzyh+xUvO7hzjVSx4im2
YU1HGEOPeDl86M/OgTZ/4Mnpavr1gGHh5IFjGjjAPgSGa+Pcq96Q1gFodwVG
Aq/MTm+DA49L+mFAfpLqh0Y9dAE6Z/1lxBXHQ0n024zIUyWArgplzGaNw2Pz
3d4m+FRB+XT26ono3Q62Rqnml0YT3wCH3mJWmK278Iivm7B9HsfhcAFMf0X/
htQIn7AMOJtjaZjESGtpHCzYTp3iQOKxIfY3lLqsmOJWHvlbg5yt+OjMqlLN
BB7IYggbU6+7NycW/ZZ1JO9lO2kX4RayFJzaq4PclKXoXpEzmzdNEJRsQL0O
bPtQD9QB3pIO/RYkG9eKe5GCZZmye9zLQ0Jb7r19CTYMLDfbmQwePveVLPfv
y7IYP3BSheSxI8aGB3fdpNTwyd0WZDK4Tywp/+6i/jDMfXNK0JPZ0nByPPxc
4cuOl9AAS5gy7rI2mSsYutLs/6MWjgjTrvu2g1PlIFBX0y08NfmQEYa5hAsL
uhzzEJQQb4yvgqEYQ5znCQQauUFl1P+nlL7MBeGvaepg+emclhqkkta3rK1N
tgmCF7Kvud1pa43QYOkae5Rpkg+rR3WCnjvGjjJGkgfUmltWvFK/RW6ACq4t
lP/0tFX4tJ0ddsFn/fa/tDiwrc+R+zVVHRI3lDnR1apmtKgX/uLKFueMTD+r
mwbvNdRbI8IlEmaC2DSC9Kz26Z2K3/ff3u2aIPaQ96wB0XTBggu+2y/k+q0u
O4gdiqC3rMxkXcX9dfHoTVlGEJRVyqHzkvLBYWwxlTzvaKN32/6JHCcrHuok
Sb19AbzTPxTQ6R2J6d5JdZF/+4AOdcW6Ckb5UHtJF7L6pJBYTWxAhPgmbKXR
Eta/KvPJwP/9oOFRQzy0kw+c/WHrAGfOL1R+9t9VMXH6tDJMDCTGBwUsZIyT
2ElRqQQFLk3zxARBpagIcV+FsMdb/Vzub7euM9OzRnW13bBabcz5rsL71E6O
B8JOPO8Av1LAswKIUQkRFWy3K+QjGbF9gGVBPODM5i2GhobIXUv+H3ds3RJM
W199q73n4OK43mfuc1spUzNUZQdOAPtEqS6S3ZAHIHdcGCcfONs/dD7PFAJD
xYY68clintSPAB4pUvubb3NfvvOpY5+nvwHV3a9mYBnoUu2Ggqr1vuGu6L7n
4DsuHZr2mNTg4BQ8J6MQ2jS+zsYrRk2Wwx/rx6pmRTYks/EBTEoDyUqVVLvC
rmjsP7CMiQlRPOflpnYfPL8DGREbrd8nxc4vkknN2UsAVocxDP6Ha6As3E3s
4XrwK07+ctyD2hHvm85zcNBcvK13ryNmskUN3Ala264QzI41zUbDZBIJvHPh
4aIVcbarDIgpup/tU6C+A7kAmOYV1NH7i/WRK/LXucb7qR3DDpNKOPsMvvtj
GpjDq6S7F4y3IdDo01PC5GsP+DOJgF2PlpHoVs2cTZl9ky9kaC/dEuKe7G1p
fiu5t+NW1/5S+X4v71m48sSkFqvltaXKaR5VjuM3q0M7xxSIUWv8W9lX8GH3
Va47f39xcY2j4TUuQVfFOcOCOEhu/WOsvS3YGoaRjgi9vy4AdgbQ7c3lNYts
/UWb6iLqVaJPas3xAzDgxcCcj9onjnfSxWcOLrJeqH9Lt65i4PiZKyEfUGcp
aoPDF5VI/yqNe7VqaKk4CYgOrKgFUr4NEfe4mgyIXxHv94zxkzKZL1XAVdyu
ZKNn6ZbqnfVnl9i6BH+jj//jPlrMR2OdD1Qr0Q7CukemkyiACo5++I6Chg1M
tAGs21Sxvc5WVPB0yC7NLyHvLPlL78hEe4R23D4dqjSoBs/Z5VjcrtXzT0tL
DKCuDfgtu3N7Mi5z3c/nk7M2RvDhgjkzIvTqaIR9h3bSNpqpfSVCajdMKZk+
ZsB/vi3EJo3Dio56UU35wIkeVOhw1e0VkFNWdAzaGCmlZEmVt5qNVy0z5vGv
DeV57He/l7KoHOU76XOVesbjVhdGNswKQAjoMwTGxtukovKUXpfpc4WwQ+Ou
fAx6wvRby9w16miKwuZB5xKd3o0YCoySkAGOlQ8YfRZLMTpUswBfYhzho4Dq
9XaWBu6DBEF8kYMX9mwrzDyIgKoSpBXzYVdyMgrszX2EBnPj07yKfWJ8i9+Z
/ouIKX4guu2Sk1JtrV+m0gdmPK7gAYtNG2Fw8PTx2/tGn3ml5pH6hl0kG+xC
YqJvzC8w9VCZVds5CK4t8HZ3ybBK0HAkTKrqkAhfXeCKTBhgUPzTl2brKGiA
k9ZELfd8C1bLHet8Ppb5sOhp47tBnUQIFPwf3HEYcvdmRVK1tBZzcd3CTWoc
voIJbkxcPRKr4Xyhc4uoUvklCj4hwi5lxZ1WyVepRAR22iXYn5PyrVMhkH7j
F3L/eR1z5vA3GpWI8SW0jTX+3Kl8AZJ8XfNi2VqKRVpLruUQHHrV93H2IgPA
G3CppxGXYXndAjscei9cBuJzXLN8iPSvRjCXU3DmNumZ5Fv8cXU3hOR75HGd
+XPGhkMMIuP3/4BToP/ttEToNX03VWpAuzCF7ohwAihDXT08XSZWpkeyINuM
EJxx+/O7pHW7miZvzMOluLmdL/8D/0Jyw1E9o8h8YDbGifw9qZ7w0mkS9ND1
FeA1SFKHvqPzaEm3iPXgllSUaEO0KqRmt+MNpNq+iVLfpmIojdennY3AghkE
prYLKP/TOCLJPk/LlGHeUynMVtP/bXmr+/wgQEz0sclklV0uQ4m+9OZk2dTr
ZCXTWrMGesESeyLHjLE3QzUXigRvoRWzma8LlXAkOdcrOa3CNngKOQv+f6fU
MJfORx3xmWWAcPTc0v1/S0sUsfn4LUfhf5YFd1gVC9Puk2ObJFe/44C3+uun
M0Ub9EgizItDHPwsZEQ69qhh1Uojl41nlNbv2ywoIt7xOe26tUiBwhkMCX68
zZOHkJaFzhwbMTJVDhEZP24qvTK1sdjt3Ye3WELAVZqUfpmm15N/cFYu6dly
gzbBDEsyQTT9GACq2iYS0Dh1dyWsGZBIX22vf5RFFQdagBhEMYBPdmwyWj4i
lxSMW8Acrt8IBzNUIpFYaXXhYwre6xT5es0Ty4NDlAjIYpxjv77JGyowTHM1
I4nSEdhcwcLFmDGHHkHZOZUD2UVNKnNdnS1qmSdGeRw355XyHKhj8kL7Z9K5
SN4o0cp5AW7MuThuqsBlZ3Q3l+ryhilGChQGKj9WPwSEYN5lEjGu0yVp3koH
EGUunagorX2qGGdSlqjziGKNQPz5zuEbZBQQi4BJJEnJHLt1w4st1V/He0v/
bmg+xrCc1cbaAEbmesQk851XK178IJ6KLmtpOn4ivQ+fqBNHCfM8q09NOvZw
N768abEO/7Esg98tEaKKD8aDEdrsRXgPTIBWhIrpzhaWA0NkgUr+IBc+rkCx
Wg0TJUGu1Mz/Hz8rjxOVik4k1TRq95MlSBSRpoljmYd2p3sl6isQ13gs9X5O
XeE8jebJTCCC7axGo3ETyMUPRU+enisxto/ShzAG1ijFCDkyqkmtVQFCFbzA
wslvbUVeDpz9drTtWDEVx/9UWhBV8al4rrlrjpl79Wudy9Sg4v2WeMOVAjMN
sLmgFbPqX2Kk4kMxdhsMpx6lWQmPQxmVh6veWS3M+Fv0WYvKtAVASs65y6sW
Fq6XHNSleTZ/t5+apbk3Z7GuuHZMyjOEYD18K7D9e4tZSADD1aGOT02X6fbQ
l9/LFsF/isBhEVo0ICUWJI7KvHx5YplB2oJm6ldvQJYa98BjBpVSb0WoW52Y
GYN3psrQvOgJ2hjiPzpTB1HVaOXB8ite/pFjh8Mnzn9yLnSmvbjzRRlxJnN1
0hPsdg2sUqgseQRZc09y4Z5sWzvu1w0usTMpPkHP4x094y2TdFqNRRQ5/ESE
TruHyG9sOccLdsv2JsDNB7oNJtfu56mvdoLfTdpQjGL0EWNReS2f9MWo5HS0
mZDk36VurAJ9XpSqER6IL3/mM66PYSgJBZ9SGIrVLQ7TwSyA3PcHtGZESKNE
Ol/Je6RA19hibQFU9SRjnNkt6pC2OGeHV1is+TD+BtsiTrj8v5gKGeIZprFj
WYu6y+JOwoXAg5+SHvvNcDZg9CwI60b8meG0PydfEZgxdodWcAkbN1PDoiYQ
C9q/mRbU+acLBFzqFCSh64Cc41kZqJbWd6RwhanAtyKJdnGD8/kn12t9uMUw
QEfLiWlbKyVyfqcqMMqDRN21AEht1lqiQo2nKckbtdJ2wv+fPQ+XFw7hLdEK
fl7jM4w2ygyzFzQl2R2pkVyT64t60s4l+zE79MW2nfwoHfEfM8N3UBi1k4qv
TcyAHmzCILYh7v+twKGWzbdh5Bulh5KLqj7hwXrPtkn/dSBwbyESHrqGqjeP
FM1qV0+qe+Ut3dv+jZ/gtIb9k5MTAfwM1APtGvZXvRgooGnkifG9ztXFqDOE
Ktrzba4Bqo51j41YwmW0e1+LeOMpTwpzgpsXDtXI1ST2JjiQI3u0LuK/abeF
zK+EFYmyO0kfi0x2bhZNrWdqQ2PTtQIdNr/QCrlEnTw4E4NShDl7LwNOiSGF
MNe4niBVOXikjk45oEQQE5AEum5gzN+3FKi78KLU6cK6JbAK6hB1/3u7bgBk
rZaqKf7U5s0RYkCPsRo/yZhmmZ28EUGogdbNlrKH2lG2Rww3np1vKVUmxSZ3
WSnLIgneC1cFPOdjgyp6aGhnDksASZ6vbumUtapWvor30sMhSH5io2bYpPKL
+uqXpU61Ig7YR93cDqEm6N96apZ5DWrpYj6rJyHS2QEOVoUUscE0SLR5UBp8
xExZ23NwvHuXiPj2FDU5On6CxA2fF9B+ABFbtlfjwQ6UfLd0uz0w9Tj5dk4R
eVAEW5/wGee1lP89MlcbPD7ot6R3pxA9WWa1nWbCoBUOtc6XVzLBUWR9S/7W
O6/dm7XdgV+/u6iIeY6r5kWL3L5JNuD1tL+AMVHlmMuVpD48HlW5qwfk9O9n
gszugLGRGyZeUon1nmo6RuTMpIDEvslvn9QRbeNPwKmso9MY6lT4JwsLjtuu
qwm+dLm5GWDknDzxyJcEoRX0d/Kb9xYcPO5ZilkAD8MW0xI6oNBTprE5wytO
QXch1YSbLX/wIt4jdoaOL/BO0tx5JlaiXv4bTdpzM7Ejv70uzZIJAkLoV4kA
V7arFL4jjEEpYgau3pbb4DmIAHAVRLop2YIT0F6NIPNOQvG3/3o6wCArrldk
mJMEvI+GPtre0y7RPYkmUc0gvgwdA7sHiKD1zqr78+NBommG2/tTPZ9J3OOX
H2HLavOpuahzvr+6LXdduOvLf39copHznb3U0UG/cfoFc4Pix5FaeMD1hJ/Q
AzlTjDZCVh2tXrNeSyW3rjTftGd/cB7+NtvHK1q5WQ7zcqMYer0SMQTXC1pG
JJPb5b14HGjG/xiL7bYQfPBFtTQs/4kbsK4WdSrtH5YJYSG8VlHBW24vEFO5
wq7qhz0AiqKFvQ1JG/N/O9aV96FEND+DSQB0FtLLDZeFUvwFolPOU1Ep9rpe
OgOxErBQYeGHjaF5Xcl2JPkOIZd02+j7ASHZ2tNMrfnZiHLkUUk4E7B7AJoL
OuZrJEylVYPLSWgw21r2DAK2jCCHvG92urKoSqZJl+0wPqGPdsLwKpRd/Yt+
8Vb+Q/MLGmztb/TjtcX9sebJIaZF85OpLHWs0ID2FM1s9hP7zztCI7+1cRLa
lyAw90zYMW3+LWPjOcc9JIBAjqIFT6VC0oYaOBjHgVM8IjhtkFj72nmLTBCu
o0vZJiLtDVbAuSqmRAc6s7hYdHVrwvSkSn1JSpgHGVBqmzIxms3hlWnOfKZY
hrP7zu0ES1TNJPr3RVEZTZxOEAYW4ld7w5VIC26O5Gf9tJqwRehEaZ7tu9wk
tlzM2l+zh9IoVaGs3RejucVvwUpo6IhB+JZ7LHlP5eoQYBy1twScT27yAdIm
4n+tteGt7Tz0qwA9Elw3ZygTn4rtCevw9qMt5ipmgHagpiCfQbinhlv8jzUS
y6N75XhIzY2ui7mxLxrstNMIvytwvNcKZgpa1ZOuvtLyTXFG7M1DGSTYAaHC
UKrWhhxBNfpBnon0yD4c/2pPRPRzBecV+Wzw9Up9zRBeENn3pvYjreOJp/8x
o9X6Jy9etyQ5vhg29oxr6qBXUC5SpyeTLLZvOFX+j8CXIpVOTA/4WKI/iuf6
RyI6+lAvCFI43yUXXS1/VVTkyx/ffkiQfMhjWCA0uXUkNOdik37j34C3H1pZ
EPMJccPOfOevG4rkfPXVShPSSy4UdU85L7UiULnD8fuBYLE3hItatQgs/JN2
9skxKCVybuERnbEo7KPMkJ2EiQr5xN93PPuL3U3aknz/GM3zJkeSkg3bVfM3
kACob1HxFJrvynt47UYgngvKGj1gdYhpyBBOTLXgW9oxt6Gwlisf5yVtgq1F
aVcspMGXdDroMTZgMTQyeB02pSYQsqyZ7gT2biAlVdqzw3ygd/k/D1M2VDfy
/NEk5s1O7gXNDYmYhUpG7hZcYQ2e53bi3kJEESQyAC5gPwzmtzPTPouDyz6R
tbnoL6JJuAWkVfhmn7IzjjTXKbLS3MFuodpZoVpCs6B4daQFXpXmnwxsJtsS
I9ZJ6uBWe+7LSv2ew5kaTQD35VIx5h6T1oshdhXDeC9B5vw9gek3H25bq+1d
/yFBcoHzeaep/guyvisZQ+D4U2w+1j6j9QHR93ORA1C15t0//9/3LspU+bng
0DJc2Q+0ERe93FzI3Daio8enU0QzbUJtWonyWCD91vKvfvQ2rUGnz2MqMkPv
apZZOeMiBDRwnEPJPei2J2B8cOagr0c+6ToiHi7P4USRnikbBvhwrO3NEHS3
bRz1oV8O8HckHjxMWdZakCAHua9slJ4jTtA9Lhl06b4WUrty90yVE/a2cWwp
y33MNPk8BEbB6xT0EtOLer1IIrhhOiZOju+avAEL158pYFuVENL9XDBqDMnH
KWcbk03b/JEZ06jl8FzIc4cnUxvKvTdbriLzvcetEqoYI3Q1+yCRn6PWR5t3
yRIAcYjOdgl0hAZPo9mfv3csModpvZrfiH1j0CeaOCsr/0D+PEHOBaQDASq3
GaT3B+l1LL+Bp0vVJpWCFmlKMmYSczWtzc8BZfaeO4ivfZJRBbBNiJQu+T8m
1BLUV7f0Z1Tj625Gpr5ELxxXVZTIUAhXXDzbYtGqE8JrzjYgKYGtGHT22NZG
VCIv/JwUl+SwjjW4mBca6ajSaqMxg11VjfhZTiyD/hdHyuPJoLp7p52hVL19
kS6naf6yaLHBe/KQ/PtC6GfkLnAUuLwIfQBMbq1NR9rMXRBdoKrMhWtarrwN
hJM0SEq37zQfA3ZICdXjqcTqdPhCHrHzpKnrttgeMQ71rlJjgCgZukaQSkxR
iVIJJSw3XL/QkN2/Kz62OEZ1NXzqqUsOD65jxo/nf20FbhB+XvWszwAikWBR
0sS3pY9Tt/hF6qhLfW61cIai0/rKEVxvSVrzPvZhZk1YKJRDsgRkaA9hxF37
T7DF2b4RUJlkMo5OhL7i/2jaERNn/ANf7JPfX/sYjvOksSVlIyaGvz+A3ALl
t4mxc3zYZeb4g1gdmTeoO0mc2EiOCy/plz5GULaiAlnwzm1xbu83hIjQ5QMJ
h1u5tbVOrbhoICU1xZqKs78hu2o3YDOGfCnckK83pMA6lTTC8HdefGAOuBa9
VDz+7d5K0NoUfYouoicu1sgAa/TyQAZ4VFwQfKSqw5r5UKhRTIqC9dD9gi7B
4wN0LjDW3SC7qh9Sj8wRGcVIIdCa8vx4MGIZ68h2wVXEPxYspele8WuOHC2L
5iqqNO1lTLFoPLO4NUY2bEVA5tNCtLnAxJTiwZNNTH5lFKAfZggs90mM13d8
4z4T7wyfEStFhyD4s0A1u8A+UiJTOpOaqMistfmyjBM8AFGQgiZLzVXiqjdw
FUfzHAro23BBSwAoIgySVOPoTNnwAlaba/AYnF4fXEAz3OiiXwtlktSm0iL3
9D4fJLAaWLvjpyHY60bbU7HqTl4zXB8gM4dntWkD7vji97P09kH09MMa1Q0Z
kx61P8+ZjtOyuuNbycq/1Bq/wknrOxsFTyTi9LAwNLUayQ0PH3Ef7QKfqAw1
KHVnaqilhTK2Wej79FvYZWgwaO3HOewKLBCyPfZQEKj/09Mhq+xVruq7P1VJ
OjKv3FZsrpZFOEVmIzOoqXOc2mupyviJxVw69nfsXtVCXPnQjcZbDcHO+gp9
xADhGxoypWmOcGjXKNDF1GnJ7y5D07Lv46mg5xKv8BOAs8V1BRxegJImt8mY
MwMwdR8GIwMtYmUhW8KHx3PedZAqNbpPxBm6xNLHemn1F1mrgS15r/qKHLVH
N60hNSCUzq9mod3fYg4lPARNxtbY1q3FjzXi1iwVXgCGTnkLiIX7YLpzZmN1
dkBo/1ekjV/PDZog/kTt6VcCSR4aUTWEN+mN70kK+CuCZv3qyhymEWpoxSS/
EvVj1FKHIICd4oGIO11go0HLX37llw0Vna3cfPvNAw4VyEyqqFiuuzmg3scQ
HyWxIlYrwvt8b0Pb6A8kWghxJxPKaotjxsXjE+V+kpMNcoFp/4tSL34lXzpm
Ba0/rHcKwqsLewngBF+2mR4ykio+2oleIEUnxznqPRazRE7Av0M+2UVjv4fx
m5B6/NHWAqHIh+thedXx1RipEoneuTSsaDF6RV2x6qKICKZY+pgiVBS5zbRI
DsI/qdTolNcCLwmRmJsC5rvJ6ASd0//yKh37f6m33yPRbk7vyy/EuE4glmQr
I+MsRexbWuxk9WofRAMGF3TzS+EOFsJ3LfW8tkc+Jctj5UJuSupAfg9YjBns
qnU0IT+WnjxpPUbFzLNkuOJphNU+DJJpKIx7K+OI2kBfxkITD4mi2K6froCy
PUjnFhHTyGL1pUv38t/kZsQz1QUjxHl/Riijh4qXEwk+JiNuRkqctfyqSprC
D2yd1CeHuk7ZJCzvNcy+rrw9mNB2UJkQNKrTs1qaDf1kgSlaIRXAnSgyzNKk
UCesQyp+6wvAT52MH9f8xvQN8GpsO8zUPVSS3eY+xYJy37xP3ovkcfISc/m5
magMvNghh9Gm5amMLSMWg3fonVN6BJnfcl9BF2fDjrIxfmt458iTEbuNuOzg
2orNT5Daql8NaZQgBQl0oo7BH8T2gOLnY5CLwiUcSQkOF3Y3MpXMUnD9ZIf5
WqEAqWrB5jumfaDOAC5ZOu/oQoFTil1tfQYbrYojmYhJE81EfEFGQYURL8/K
xdI9npEfSKxafnWvfw68f2uZHshiR579D0hDn7h6YufaTAa/pXzhAjmvdrFp
KzazubdpGXibuD7UpnKaUiiSEWiid9h5r96/HE6+dpXSZn4oisAnGKKaPmVf
LRTD0O3WldHoX9GMUUooV0atR/h/AKxi/yGPNNVUhC9d3YS05joYxzEhaiQn
LWyFKgkb6bfjzzBAQ/Gr9vhvvfH/UEJYzkNpTE4MkDz9a1KzgZOPJ6FkuYHd
mV/Xyy8oIJPeraG82ZDhyjuNs+u9xIw49iDXZuqcubOgCTdUEGkJIVuZrSrP
Y2rTraGvtusnqtvB8FS4CgUkvqGKxXSqbP1PM6mzEsTQTOwFITwkHgaMXZ4E
Ul8NbmyFxyIftT3YLvk8C0kuQo/c9FzxWJygtJLOPDu4bHzr5aWKAjbZ3EHN
tMeLq6VrXs2ll36oLSS1LKcQUy883HzBKH5hpWrqrkw38JGwwX1rmdEsMDAU
zneyX2e65Y3qqRKKZB0Ehezcv1VL/hwXW9S/5XflEstIz5yPoMMby3C8MuHN
Hnff9ewgofVheeGtjMMvrBPJLWmKzYgfC1Exm2HmDAgMlfcdTfNHcJYg5CkY
qUGzeijVtp9A5H9drRkT9XJrZzvCoecuqTOVcxk8aRebeqfNU3e2kWe/mmD4
RooQFXoOlol01Hwmnfh3GnbELrF6dGXxddpYKsIkmpM4x8+oRZJR5uXLYYtC
gpOMJq7RBVMi09C9N7GbZH7gUao7nPHUbJ5AkD44Z18EhWjxdJNck7GyGjAu
HuwQDNbMp/OzfqcFJiF/uDzaar2nNzJs1UOdbFkuJ2DUXjDL6HrlYqiD4UuV
ElPVl4fd7Ie+fR4RMK1aWkLik1MmA+/PjiUt30TzReG2iuKvzl5AqtoQa9jc
cl3CQl5vcq5Wj7Z8DVGu0YQJX4RVEUwjda/bwM7cSH5297/w9G3MPa83L/GR
u1VCs4cBbVyk/BzPFh9DorDtvF6L9sLatWXRD+6BWrbA9AilOBhD2fxxKnnl
5OZJaBhJB1Bl2T63QsJvj3Vfjmm35NX1VBUJi39OJBKmly/5jyN7xsaA50UO
mzU2tq+wlT2fs04NvbJSy3mPUqg82znx9ju1DWHNYVsfNwO9FGpSNZD51z+u
3Df06C65fszy2b8ZBGXaKWQ4D974dwpkwNAkjajCE+yg7RE4EVfNjQXPJSQj
hvfUSR1pcG0GAM6op+Y2gU3/jfn0fFVWMpEqkMx9amD8iFXLivDyJ5Rgoiid
BQpegod+y94TMCO0vwBXQjtCZWgL0omz1Wiwgf9dJgVtwQgpkaOGWJvTbH48
EwDOOW33vdk8rPldCZVDs09dSpiNIGoaoQdIHUETo7k8QILvs3hxAds4YbzJ
QnK6Lx0FdBExV17mYhfbua9hFwbfSlF97l1v8UJ8munbhVJCP9du7hgzQtrC
uk+mw322IsfZEGDJ4SSvoYmkYMPvUoIVI4b5Ix/Tr7KdWGh/Df20Hzni+V2T
3Xgo93nfAsr/Auv8zp3f1qQQMs0kfoRC+T5CeSSK60+JftbO8VGDvUSbIzaw
VDoSstNp52wSoSdXrBr+VXERjCZe9X9Wdk0ZLeYyZsLS8rdT6tWOsemoAVkF
bEKzmBJy5OtdUGao0IzW2aIjvIte+KFhbBk5iUHd6P5UUwiKF4QwoMw1mvYd
06QXNlyMrGIGdUze2z90H9LOpAzzer1KUCuBIChhv7bUOR/5KUe/+7eug1r2
jqpNiqNu9aKqHhNDp7wOt9aF6QPn7wKcXb84hJhwemru9loiNKk7J+WjVYX0
nmiPbQDdXERUHjjyEOYM4FWdzABlOhMt/43E8fiLifD816ktG562x/9YTbZp
S3qzB4pNEAKo5L3EOaIWaJjYE4bIM3eUAc45VbX7a41vo5bzQDxYuS6yu45Y
xcBqKkUfwzwRYKLMb5hwvBeL1Q5tkXoBQr8daYhpPDdvnR53hsCtq9dscP0Y
2JcxBqnmDguB0Dvd17QkuRCbe93+25bodMjs7fKncfiIcv2PZmlr8rxaZ6t2
mzo3TpMDOm1PC+71c2kmrk+RG/E77R6w+E1+BtEkngOHr2w6hnYtNZLld1ck
s/36swQ/6gQoc74n+uPP3ISEKgbIIKScU3bjUuPCXHKLyA6knkkd3BtVuU71
8/93LWeb/2PN2yJ3azr3RyBUDFBBevTM2AKmER+3jRuFYBi1D60/W4kSetPG
Sz/i5bF08r0QyprXi9HY8YLuN3YhXTPKFqUU1cAsaHWN1J5ODgRHU2btXbUs
YPjIyAWIpaXp8sJWMZJZbEhjlUC22jPyMBcSyVffYvoEqVXsZNBi+WX6OMSK
wfKZZU4Y3j6tjwZnjGZ+Wq8t4X2lTMwPXhHcz4IMRRL4oAdOJw3Io75QNa4e
Sfbq3PGSYfxHhRuOuJtCXyPMul7cfq1Cdf///7maVEDWvp3NqTCPGgMQM3Fn
uWPBoS07ievaVi0kgnQYzdSKvPajflo7RpTM7e29LSer4aqhcnf2J1xXyxPJ
674AUTongYsPWf5L+dC8Jgu9cSxh06xzv0a1pTgI/XSLYxJrCwyUdR60zHWH
QGYkYng8a2jrlltBuP1fe4e9jaWTsonBByAXl2Hy3FsyZ+b/EcKbSwF4XnMB
8cFs2+bn4kKDRTOP1qAw+kaSWuPPKfxgbbpR9hClgVA9/yKwk5suhO4rRv9U
lV4BNsjDH9QyRMvyxITEDod+53uQGoQeEY6tvuB2PcEJMX2AjFe7cUbMe+g7
Czsc46mpnWqsjlqAuRh4ok4/7vgKIYpIpMwOWruNpeK8tTcitF7b8CPJvoJM
+cLCeoJyQiEwaLTWI6jkOtcA0+8pz6LD1Tz9391yDUbNd7xFIez8AsqN+lCY
A3rhczL4/nnP7Y9ageCV2wopkim5dDZrrv+4IIKCy5+hOfpFvGXINOoO954f
Qjvyi+P2XfqAXvUFmMo4foqQAQmeigacXA2n6A69Dh8J4etxsl94nZ7GxM8a
hEndy7cjxGDAw6FHp1RtQA97yuDUQplja7TZOexM+IBlw6qJYF7lfL5uDD1j
EPWULdBtfbfciilU7o2wPrTHyEMCggLtccrcqzpcIq1lFvaJIOUknmUNE3ZJ
9h73tdw1xRtQxRLs1NrpHdYRgfbTZQTm/mC9ckp+SjRvdY/MWwBUUYMLPInS
QHnVRT5f0V9vyMURyIjwb+44QEXts59D2qu2Z81DOP/uWp5TG6tiKYRtzy+5
IknEh7ayToXcoVI3xGM99aGEtNzran/x32Cn7G8eLYnjDH/yj3teaZpqXiO7
e9B6qeaomwWK3Kz8SWnJg0+0arCwfZVQ5QLPSp6BAyHZvFyk2Hx7qpplwvFa
/GfZJABp56/o1jLC71O9Q+z5GGvR66LSI45fdPEUHCxFjsbte0V5b4A3WXZQ
cPjYQ/v69mRBKJsBmJCRWJGAJI+ipNbOeDYlyFFXmFNtbg3FsJ2reVgNJ8kw
XESnMaJ0NT38vBP7h4UptKJB0lXycJIxSHjqxBATERjD3kkqYdJvEh7Uc/wg
HrdaMdrrYY5glBJhMlkM6Goz/SgINvPJ8evJOUv3evc2aXu9o0Vb1eN1ik2t
EBsV0LAmj55o0rpCYTUH88fspcmVir9iH9Sf7ASUMe8WZTS12BGGh6hYA0r+
iI0qOAhtBbdjgP905Bgix0NKEnlkF/gak03bVWOyGkIm0RbgOZjiPfYa5puI
0/j00G9RUxa/rojiTHCYp4fSnws508BsAhcbnGfG+f7LWPm7RGk/lbB1oHbz
Z11OeFsBi/r24sWAFDc65+hWLYcu+iJ+3Ig+HRSzP1Rfk8LkT94uJRND9xnk
UCiy1z3LPxiLYNe8oGQ37h6wxzpX61Qf7C+7x2c8T5UyxHXFD2rfCwLFqa4s
TWStHcp6FYTqvxV1Xb+etHyLYwg0rxkg0kbHXogBFyCDwUFqoedzn/8CSZTR
nVNtSVkiFv7xiI2a6lpyjU9THSNv2OxaPML83/RMELbKSVMZ41lMFMxB+hQd
IJwusXQMkZmx8yri4odThAvubF/lzzSfgRR071Alq5d3qeAGw9H9PWd5wZPK
BDGwLE/nRVbjfqhYxVrDJZiRwfeaDu0Y5LpTtJTpU31UawSskx8rBoseVuxv
oB7jM3/ZzfC+0VkZrK2hW6pKajC4y5JLMHT9ryYnGVSsE6DyFX5MoLUjwcMq
8bPDwYBmM4zC07fczbDLpfKBbGjSHldy5sOInnXdMCwrzJH9iBHU83blTyKH
j9vDObzTuK8uY9vxtXFuFbfJb8YBQr6vb5KnTDhL0v4G2Kf1C3+7EK7PLOPB
FdV6dssgnjdh3YYF5Ri7DF295klJ5841QKBtO77fW9t41P5udYYuGy6MxWCY
2OkVGMyzft7U37Eh+HEDFWf+CLn49XzzFDjA7PSleleoQUcO5PTyrH4UC8FW
3O2LXDAL+DzEFiZPS1NOU5qrxr8IrYyzG6e9mbLbUmyfv/pRBuir+astVe3c
n7/qszJcbOR5oZOZ8LkxRQs0dlFgHiH7Vmexj4mafWiXpCmSKjAWhOirQCm2
ANL+Iouaoc25HS6AR/s2U6lNivD3xjoTxkBqWwNMYXz9jy36YUZH0nw/iThI
CPaFn61IDx/M3bVc4vNgvOvcjiax8stMtObgKYl/r34Ro2V5vmyE1MsV/uY5
iSJug1yqbsOSDP9gHzJKYOHEVfpjuUXGJF7A7yl4sJPz1m5Wro/ltC1qjUt9
o25G5Zs8QGp9yL8LZHt1I0QYBBuX4PPmO94d/ibeIlZKUxPs9vmKXPHcvtWt
sHe1NMA3P/7FBVbe00f0zqT9V8urDg99Di47vhUkqBOsHANTqUUQpWs1zThl
OMGqvFdzsKAcoaUMhWyYurQV5ez+uiuYkEBDNoRVkSJhv0lLB5PkNt5Lhs4C
KIYoBna0tgEUvdYAI0jnXDXyWH0tqHBaDCFZXBvQB9wxBoqmwiiW8nWXiXHG
wchn+bNtUmm2yKXkNwJfnrk6Y2bZ9mh8BbRJBXidNL4p3NKPC097p/NMZgX1
lGpAtjBAH85rb03aSuJ4ppGL6yy+Xwz2H1GdTwtlbNAopchsz8Tc5R70Ye/b
LKqXvnIOYqpKrFx//bswXq1gvyPtDoe42ThaEHDUpjbWD0lB4xeqP+FNL3Th
EZUQ0EWKKTCUQEfp+5fh+0wLvDSqDOMe8hkzB+CDZl+ZeCoVsgW+vt3mmVjD
dsRZGzJ+6SUXmFGjpgvrT7cKa9MRhIAp9loKbI/nSETKFDx8KxZtsaa/OuAv
GGgwlk4HQi3CSfVrFhFHVAgwD+g5VnpB77v6tqZ2m2H7xZ8NaJx7TdHtJw2r
QMqXghB7zDpaNAMDywONzBgwpblD/lcoTdUI4TqyTdPgmqB1hgeWqBGiwpwa
l0iOmrhNjyJvo7Qw5GxUx5wsxsfJb76E8jVi2yC++xymvaX1xN8qJYKiVfOO
9rSSvay4cbLO1FDLteN3io3P7aGdPCe1Znfp0/aMiSBOZuNJUPCHXoyw9Q39
bgFzGnq1Os2PMR21DAZGNkOYz6SvWFlmtbitLS+Q3KZlu0EKz0/wbUJYzUn5
AFgCCOLyKkxpEwPtTIaCAPm2wj03BiuiEVN8yxEW202qAfRy23dOLH9C2bAr
xvuSGYDUmd5qUMS6MK6lykN0txIyU2EO6x3Xii+cVjN+ioLz9pcrGps+QyQM
x5d2zgWRFF7LaLK0VFvnLKr5tUr8AY2zwcvNQ7N/ajORUdVRGUjgWvL/6M0M
coXKkqShLFuaEEpY4cHKDqK+1Ea6PzfW3vYoC1j4/2UtaSdJaROt9VTDS98v
wWkOqT39W1IUbk2kHLdszpaWyinQMowuFfIZcx8M+LjfGehGD5ZRpeVFHUHL
2MwYCe5khSJZTqY5rls+9M1ei01m52O8/IGi9zb4Ng+db9IcLZGMAgBvfqBu
czzPbc5g+eXOZVKpBwhjXkEx1clw+uGpwJsNk6mPBONOT1RUEVjIPJAm2cv7
Ai4FQa6cZV3QTRgxep9BzlG8pLU09N2OmTIxQG6aoav5iqzFPAZgHbF10uR+
sA4rE9HQ+yZsWTd+bnMNi9Bi6DWOmbb4Ix6pyj7YUynKkj/LSBwYs7fQiWAQ
lPFwIhne4t+0ptRTomz8uP3sLBdznAiX5PCggejICSbnRj0nQvpFMRzapGpA
CD+AdG4wJS8+IFdVGivo+EY9CJ1RFOzNgNOtwfKoAIPOPZ3bc+wm4rsAIpKV
VtfyA5I59N+EoQAsEGSHW5PP+4XvvF9ATUvKvKfyP7EOGkEo23zjloDSMs1h
SYY2s/2dk6H2usDS21LOPe+xzAYCqwwWZxrxWZdrufLEOn0x/p/SSMHdkkTT
EO+YsvnvPMq64DRi1CfXhEnf8zQcpT03xKzVtaw50qISUu8QkBkYI3VHFa1p
ofdSxMbU6p4WkFn0USSH/870RJoJqisk+Kkw+SxUuKgeA4+t3usSxsBY0CM1
gdBPmcx2qnzd8NEEDN90uZwDofemL5IXOG6avbcJSE6sYCI+mSaCwShPA9VY
1JzfTXOvl+DmZjOsm0Fdu7JfrEHIEiuB43n1sRRHW+xRNyF4AoHPO3IyLMiD
lQ9L1qM99oJlFZeKxAivCVEX7fO9vOBxgO0DPM+2Hc+feBmL8s8sdw79EFNd
lSQaLedLNwsjXn9Dj8GMYFANR1HHxKYUscJMSndxWWHKidk/d6moK/0u6rDq
YO3WkxJnEe4NXAuwIyZgw0kaeH+AnDSWwTKl1mvmKw1k3aOKNUOfIkJp7t/a
LjoLASK7Ye40jBUDyPY1SC8Ik9CqoaZNh1EWpfIArKgLa6xoAbpH19kGfaaV
tr6HzWcvHhz5BO6LfDPTRwR3dAv4rizd/uiAsD39i4FSKazr9inK7unAZ/OO
1HSmPAYjrsA7rgIjH397eB6t308ob4P46FhJmaopB0UEOPIHWUoH0F+GXlUT
MX2BvN0uYBrBgaNMVFgi8Ptee/zuFetdzaxF5NC3erFWFlgLQuRDsaAfKE8Z
JTUG7mXIAStgUWDFxOSnri4O3POhrcYFCVPuOSmywOfcRcUxdYqeTl5RQSrj
HVtzbAdmzOOKcyn9dUTohuBoooNA6ohGi6QXXFqQ/Ie54YKrgSRI3bJdxy1q
iIYHZFJio2gpMu+0UguRF2BbIVI4fwl+eJWRZ3ia12NB+Jm4zIxIDyL9O6KS
KSbx7g27YauCyvT5vrL8/QMGNEg154pRPHt38e9932fP70wj0bSXXIPIWnyi
0E2U3k8vsA2pBezGnHTspSM0+7pkSOFO5gEDX+GSsGf7NW/p3Gm3+fMd7h4F
WryP+uf5ZKXijyLLBb0KM4GpmUeCBXtqaoSH6Kvm/StcVNje5YE1LSbaKnMb
Sj0cx3QqzXBLQiDSkgmhV6TiA0DkllQjIU6CdDec4+vxJueSCgGMcyWZGiXX
rNusDl9bWwJWzfxWf9ziyBwG1InAj1qzRHmRPUMjt1QXX/lBKYb6rmTy2R0c
m2rFK84YZtV/+2DE7mGMqK0cTqsoD7Pjc56TE25E+p3gpbLCbaPUfBfRQO6n
mEg2g6rt4ENRJrSkOi2RWNjLU/2v8jsb42OgI5ApyT9UYupckfEslCXI/XJy
MAAfhpCdWvqexr1i9ZrjWdACu6gXZ8IBoUq/DapHI1+2qUXF/jXVxlLc/vBf
Fu4unRGsGOC8SKSqd7pjwFVyWVxkuqcY+uX64te8m4cy7C5ARR1rbp8s+8Rp
mwJhssH0EbH4d+y2aND5qWtQsQ/sfvg2+CUD0t7SDtZzb0eIbg9AzU5GkuJ8
Z3EisRbcisn4HW6Hv7gjo0ZrnR8hbZJxwQT66IGxYKrNuKdSDWqFV/X7FP3q
ffLE9uiJF04W8eO2tOJxFL49azFR+fhONSeaDYxCC4TAWL6BQ8qf5+m9VZfz
bcRpM631c49WyXjPETdf6m8RKmS7sSzZR+c+NWDsVIfG4XKNGjb3yWU9xZJO
CNHsCU5LGA6u6w03E9rRG8LE1OfrhPqlW5sS5RLi6R5GJdIkufMuKBisctB7
a7OQBOz5LwLI+QZgiqLOq68wSdiPVpK+IFb2aDVLNPKbkQtmkXGbbbmSlyYC
aFGUdNYyD/aemVt+HtveBqxl/90mPUu7Yfd5JrRjC3m7gDUkBPNFm6GGGXnU
uWVHYxYJbdTAPW1hDraZq/aTHfynXESwSQ33oofR0Pt6vmsuYNrmqeK9oVJ+
Lo0dDKBIL6+DTvTP91yhgkn+aU7oGnogeuVLT5FvscM8K15+/xUIu3bEWEJa
Ggz5mLDqJeizA27A/A9roOVE9GYh3t4zomr/Sj+MMi4vz8Zo16N0AvwuErVc
tufRZeSzMZteyEhvTfezcONAMKaYZ4WWlysA+9tah5joxt82Acndbcw1r6e0
GveMM98TALTs5A/zD2OF9VckMGC/svx/M69/JxFHhoMpOChxE4g4MlJvg0Yz
8ODGQu1+ci/DEfWb2zw57Jv9U4zdOBUuf5Be3eDz0tAhTIu8FjXl3dJW9aY4
hqxqYFposPzhMM5woXKMBcPy8SM7uDadWSsKCJ+BjM4FJouhjhFV3kdQr61/
NQm5mhfSLhaRV7k+7kzvMZMESV6y0UjbsXd41PJg21jbNvVrwMC0PB63uVeG
3gFtuhRRwgndFfPq20F1kOf2xCtesu/57QGWmqrmu40tCipGsgxexXdEL4Zn
DAQZLbBXGChJ4gqLyUJXMKvkjlNqI1DxPT0X8CV8GU/KautFtt7FrBHgfCk3
MnpZMyBKFpqYhvRgc3qKXCTV6qqj0OnbXfZpEF9O0vI/QxX0uP2c84CTsn67
0HqREmlekjoLZMOxegYtRSw4eDiXq1MBQ5pAULRNZ3REtuj/uIrCPiZWCdWk
H+DNqbWWBCwMTh1Ca1LJL2iKyF0ZLZd5XwMvTtLxJL05NLC8fyuG48DYBAox
dydxYaY/KMke4iGYoWKiybRqBTp9PFKhNEFhgTTCHL9I3egNmxOQYmtDRa97
e6ntOUoliO+vgN5o12XbhYfGX+nDbj2Wc51SUF5EGIufG8cCF7XiHedua+/6
lpCRk+gKxrSAYXWOddwItxGpSnYRo5sp9UU2Mbmq4gttP4LTpGrM/HE+gLvo
ELrYfo5ywQxVdh6KqJWiB0CWWho9PMD7Jn3MRxV8idKBA9II51g9MuutR7sh
y1xP10ow5qf155GL8fOyDaHy7ZhaLkwsY8qvD25zSE9CG0vPnyuB3s0kZEPv
DmeSedoNKU28Mz5DUo2Rma4UwkloBt9ZD1RZowajxk4GYmQm/2+k5CM6fant
LGTtsxAh7imW0l4XfV8ah02itwrmnIKE47h74yke8yhHsXsD+jfaU8+brdX5
zRhqzprRuNGb2cocIdcKWFib3/7/Popco8UgY4KVmPEAmessqitrU9G0epSp
EHcpkR008/WAOPK07ShsvkthCcZ8R/iSElc6Wqoyv78eONlkTAGphmTdMff1
Bv4S0UUlv+3GTgTtb5qvk1DquK5TdEvXp8txhIKUBwZQvabyAj3zjQvYt3tG
Dj/wcAB27GwR1xDFh0uWPYg7UHOHxex1yyK6CZ0L1g0emfHaN/EMDI3KKybw
uU++jS3DeUCF+0j4AkJCkM63I6WMUY37URzx6MCUaAWq86yxUINSZhC7KHdN
GHeMW2AMgOq7f7P3qNC627gUbxZOps9OO6V4otYga//VjiE0mspPtKTqxMh9
uXbTbdrP0GX/J9rTOeTu6klZw2WrY7c9XqQP1RFV6ioy0x1BjjuhM+KbnwHH
jOeyrPn0chgKl19U/Ib2WjyI9znUx70TefeOxe/4Wqz9WJR5SVpXX+djKPwW
v1UPaXzGLDF5dKT2oWm5PkUpS1cMPkty0iXcn165nABdTGwUIGEUU86L2wmG
beELxwOGMFhOweO83eLb+HOzS2fnAp7taO63OkzmWD6Lxkd3LZry5dxsOmic
DkPqyDOSPgKsD6FrWhpxyU8m4tf+Xvl6IY8Hg2AEyypy3+94A1HRjVPFP58z
aLhMb1XL9X8zKiYWNkA6YNtLO9/f9I6/3dCzkFCDnGDMWXKE5QI71a/gPyv0
hCCkqLaGmOnpypH0XrK/qUmQ9fJbAiP42eXOOTtoMn0mw64R68HFbOz5Bikr
Vt66gOhtb9gQr6a+UwsI8d7rSFmFcWsBqrHM3+eHvfYwZE9zkEbM7fMM9iIs
ozRY3b9GJodxcErPqWQOQL1HIvHsqQZfPyCM6F8dMKDujWjY08/ReFnoVomB
jsg1I7GwwqwACc8IZ9xTSPwJUSWP7Rkb7GSmGP3QPXuyUlY8fdwQFq8BuT5L
a3qkhQOU9rFh6f8Ezoq8ZThhIOjgjdBZ78WIXMiQWObsIhZoDaOKCn29kLfn
3gQw9STmS4KhCkvZYM/XgCEPfDT3fWX5ygaCUzQzjPg1NOQmmFBiR0bKCEoq
RfMha/PUFVDkSryVuvDrsEe/kPE/FmU7ee9ISAtBmLXdX6pCSXH5IUCBvsQe
3uf8m1Pwj/Em7z9EK5RBINO5yUDzMRq0L+ix0rpAA7FTRDFYIixDUQeGG10e
Tm9A5oyMMgFF37V4Fs/bwSzUiuQ0Lqly0VNfjoqWYc5rW7Vbm183J8rmH+L8
CyXa0+NrXRfS41TxdgIuKZFz2DaDe6N0/UQ92/Njcw3NY3qU4Ht9b832Oqbx
KAyUTCqWTi/uIBxA1iR2RwuQ+Wbdy3dXAFsJgHejBqCt73CpTYptQ23OyubW
4ayDwIn12bV3pUJk4Zp3W1scX+FzMZ8mtJmwEkj34dB0vVQGKhjVa25aWdNd
mIHWQ9Hxy64ureO2+WIfa4JYxSEwyw7auExLgCY2xM2VzJi+DEPKQZTgT3GM
IYdfE4wICsda8oYbGnE0t74PV2mb1zj9ujE4bN6gN/0z89Omu6OEoPWHd2VW
aRrGR9zoSgGCnYy8Y0Nh3E4uwNO0AsAU557aj/ulPR2ZlTciGk/D+Iu7HhDn
oWcP5n6zhkGDYCnhHm/yqj+qp6fcYA6ER8aEcvLFCWQp8AZCOGfkgACz6ZG2
bIHs2/C8ehA4Hbxw3/PYkHjCkpeUQwEzjsevTZn4e7GH98HnTzV+3eFp0rV5
zmWJ+coUp1Q28GLSVzCEsAL44jGwClFh6FWQcMySasAEo5w3juK3wWWbbWgu
1/nOKd3DXOB7JWiHQGHRR7s5W/uXyUXXMB5nLEF8i4Sthpbs7fniLHlCI7Bw
6FP1vWm9FFDNcJC1QuRoTe7rvnfJgbmdd6h/fXwFZrO747oc9pNUTaaqpIqh
DqZz88rLlw50mF308lHk7idVwVAiiJ7GCaNQVwQGB535H3OEZZxD1E5uUSt4
NxABZd0CzhKlODLelhfAAFfHABvcBREiLl7F0+AM4Mu8vDp2yV6ybXMxXUSa
WH7qIbQRTOG1lxkm3WuyaWR1pbDGCdws5jdS/lu41ZHd0Y7H/QgOxtTDNcUZ
AMp7x/wNErFYQ6W8jVo+7xOQezrjNqZweUEeVGcjuONJoFIrrDVDUzBo51Im
ji4PeQkkIYjJau/2gf/Ep2Dm2U/zXBkXY6Eljs2ryfMgljx9ZrLDScffb68y
/xMGerHykBiBGNcIrWGUmWbg7u1SalPllgohmvy3QHzdowVbRozTAQX1WMbs
ekUxAX9HVAQGDdWGyC1wlHQIC7DGegoHMktyDFBj6wfMZv5E7rb2cK7mqu55
h5ax97vLdHy9w3h4HfQl0D1A6n4Uzbm0AVnuxJyT8Y7lhrCMGmsPRk/OUODz
LYgM+vU3oOewrX4cOdT5KA0wI28Iye9hEUawOcXoc3hTejH7I5IZoV1R0Aap
9ECR+8U3d6nzS4mmnmrJ2pJx6xaZFZsb/Mt2+UMMTflCLUhTxfz7IfuqDsn3
hWQxAd510qL3YEP+syJt7hUp+a6ZXcpKo1uwz+ZhiXsOKWBjKTEjmF/nQinH
tEZ1JzXbB9DkbKHpSnKwA7HnQ+txGZie9DT5JK3s+cabqumxBZyqe9+zKbEN
LGkrZbo4zb/5f+DKQasW06uWQQi0tyWeKoIqTjw7I34pSD/c9W2+ltIFVdCK
Me998xdd8+U8wSub88Nc25nyUMgeossftkqaRfVkN1fIfnXCqTwvqSlJtnnL
jdqtsJ/RACdDTm8D+1DfJDpilCVp2rOKPd0H563kA7whh2x7GA3HYZuWRSZy
ICe0/YwsJwyxux6+HIpvVYKJJkfYbjUrIOshJJvzu8+Gll2QQPdQTjU9i5hU
zMT9sXcFcIw1ayi9RS53N+BxVJJvrhvGAfyJovNRd30HxxJsayiB+nnCBOWG
PtPeTgUp8HQVvRd5rvLBqymHWwtagI2U5JWiI2NpuDYHx+Vlp3GBRvNEIlGK
+2qH28zzxvhASljtElzmftVFr4atNos9AnZMq29Y5M227znkgRJxERCWtrPe
zjnZCq+qR+z2+h88ywo2j/w8MFL9cx3XDJzuMhiBXqOxEovyi+8A+jnR+UNC
Z5EZOF4hfosAzn+1klXxi1SJPzSEfozMlAADEohK5aHBx4GvybFEpayIRhqq
4GNPo5v2ywxK7EsUtSpGeAYubCLbhy/5P6h7iCFCalwmM0YH8iszR9fuJHPf
T4Vs3RbjM9ZuNsnvHSYYq+gbwm6N69SR12H/ZnD38C2uvdnGFYMvNndThB1f
FHVayYD2pl9xN9BOgYOcQ4+eq8RvcWaZzrqwY3+vh377noNyXkouGoKqocrD
WurMeWgGR6E27OYbngRdPYuzVVq+AMFkhXaVZ0eWpR2ukUpXCm/EnEtqqO31
KqNLFNXSqL9Or+sH+cIDBMIiSuhfIIN8V9nMBvLApbdO0IGXdZ7N6vVdpVYz
gHq0DpoeWJZWgYW/XwnkrS4yrkUI5+hFQw76I1UCAgSrwi4kLrM0JK7Zb1M9
KKXBxF/2KIuaDb1i9bV1AsjDKtxdAsM/rM+ATqbANQB7fbN9Fps7Uo56BX4c
/TmJugPc7uh6LfDc4s/VUXNgz2Y8K76UGvxtk974/fqe9FkkeBQ7WDI2kozO
nPdA7oEUnONCJDAMHzk3nkeU9gb+XUVKmrL/Qi5eURppkUWq+6vFibrSEYGR
exKclcJO/j+CyaTOsevWrdY6j1OLHB9FEHwZcINhv7D+pEyiJL1r2BoxaeVD
FNd4Oz2tVYAh0/Q+7mxVuJyBbiF2wIcBC76S+uqr5kjNho2M+JLJ5x34AYFp
DwWXPThw5Y3ZcwzIkDcNZhDjs1khRHsP6db5b78HZk0SxbvU04OYUOefX5ka
gjtYXYV4kvz+cRNriJEy+eW9fa9LdQC1JTogNiKsdU5TZ405idcWxP++7l5U
7gYnNRgFGQMd4iZpn8q3MjOzgpS70wmeyXLWiuRfW0qU9e/hGyp5yWajihnc
PUXg9UkSKJtUSSjInX79i0muCJeC7xSAcLUMTSEqzAwzUFqgDAhPuGL1QhDh
K4KLQT5hjgB05EG3YmFQIN33feYIgniYZIjuEf0Z/16CX8kapAsmGurJtP8W
Ou1nJiXJlgClSk1Izlw2/klcmv9Pp9hYG/xbHRK/K5CJTG4bHtCDsLW83Z8i
w8wjwEHS4J3JPYeSOtjLidiIGiBXSVGu60xnu0M5ED3LHNehjyOafmjbm1St
KBtRn5GiVd2+l//ALAqea/T5M81xt9Qj+EO/kjn/d2D4j5wpvmmH/8Pbzlur
6qi3BMPHBKTWHTi7l5C7r2qL0cJlQ4gJJbuDXZHem/YEOhiYeQcWqzUTone/
74sf3mh9cxhBj9NoVNn85DJuzKpVHYK4+s0rV79ze9TJpGH8vmatwvV4mpOK
0wDE8C4o92c8/EqycVy5jrT/C7e92n456w3T+Jz5UtFEvPDObtlrCZ2NKLMh
EGQ2JLQPTaK9HCNQY4bmfW2Moz94PNFd1Pwm0Zx3+72NGVEkB+qZhCGnM6Mu
lgcdRu17nV+Z1Qy04ykFotZHTL23cH+OlDcKqr4zsGTy8LuofgslD0NA6sq+
YSFtvRQdoXwdNR3lbUq0wAH3yEpkaMnJ59haGZcQ6mKopIsRsKAAaSr+LS0O
uIK+oQoN4kVpBWnkQ3M16DAQdBMqoOz5zgWEBO/vovD8dLQ4I4ZxWv/OS6Ef
XslG8T+8+KwP6CfBAsT8XuciW6l3RrntKbdV/70IX++fLMjU5eXG7Wqap3I2
1ktblF4QwLIpeRaZGtvJJP5pq8VP/yIutdmiVPiVcfJxRlmtjBdTlQWnEp6K
/oyykMmbdDzRaK1T5IeoXTr89atP171e6rdk2kquF+EklmPRqunu60SwKl6N
16acEA/dMHhrmVZnazEJnONOd3NVSZMXPFnX1qTzW6tPLkPmqZM6kr+5Zql0
21LRPkN1FxD/CUks/lh1kOhU1tKEW3lKHibnfYbj/jAJrNu01eNKMz+2fcms
RZyyAjuUULKcauw6lYcg4E9FHj/lFmCCVIJDzsREUl+DV7J3YwpdhsY57alp
EONf2XDUHkEscigi9PaZMbhNBHt7IfrJqWzlljzlOWNO7bpyMMhVvX4M3Tl+
aV5QLsRdA0VfWBD8EI5SkTExqr81nKUEa6kdXPaeHdZiP1Ik5+YSFMOMiT94
zdWlSBDhCEby71HQdG0yTXGThjFCGPOg9yPrzityJtfxa54S7sQBmefnAyfm
eFxYAGiJUCNuoUIGC+GSyt/wSBaXGBu5TOUK5Zsd8twr+zHxmNEeteEk5w+k
hv0Iu1Wd3KK5M8ylYYBWuBa7zoywSKxFmY8vvKgk+J/SsM+1YrnVfp+CK9vo
ePfT6rXC+0I1unJvGrjaVjXPVMFj6rZdXyh0npOVD+f/+Alo/WIwdQBA9MQk
arI7lFOdtj36O7JRi7KlBcV4acfGRC/D+BVFCSBnARx1qfeiV47fZhF57rFJ
UZbMP7LlShatl0tmcsmS19QO60lDH2X0q+DK8ppiNjhW6AJPJoPDvBd4TMNb
cYQ5RuzA417A2vC0QuH+HwSEiYpRWULvIMyirbmRPAueSEn3j3Jz90sHwRMh
Q1hmhSHDaxvEy30uPGDtQXtG92xkUrePsH2YC2vpWfEV9Avo3sP7GBJJfpNN
35YSq9yq7JI5U624i7+v3nWOw4wc7dDc5xKbSFiH0z0UNOFqxA0FAwN+eSkL
mviwM52vjmO1DW4fiuL52qihiw6ZOgMbC1FOrmptf23zh4ZDvDf0SkFc3xca
tiwM381glxliZ4I3dr5RLxxGBRXHWTp+/F2XfIPAqE+P5eEaX66TVCH3YaT7
oH/zsIaV3QLNCVvyBuKJ6gsGhCX7gWVQsV9fIcnVl7079OetuG24eO1JF3za
2mlAf4/XswdBcbC+rj1W5fNXH2gdaks+UF3vlE3PV514LcSX5X+u7R4BOhb5
Ln4ac150mzeoHIP5PmlQISjaFJU3027Ahhfu4cLCADpJsPi5oFqXWUUnmS9k
g/oG/2h0TwNc+b1Q+b1D8uTgNGCnTumSugaNtlYjhwvxoAfu4uYtvMHPquFw
SgYvGzQxV3gW6G2l65KivGwJmURlHeIUh40eS16xNQJN7jYakQnUUrp1xf7m
0/TB6jLF6K1GLL8ypbhJ5CRc1MgjmeS5PX7O+Yy8hlncdqj/P//WIaUxpcVB
HMw9etPjo7gYECTx89odgcrnMF9ttbqePJDYFkkLWJLlvS/0TjXh1dF5e0Nx
8NZ6YubWXNEFBzE+ABW4o2xa39ij632nMWjAVJwZBC8eFnCQyVHKGg9KZyHc
mL/Hq9Jn6Mw3HaBZ/wq/itIOWMjemc/RfTTh3GfdQWUfZvAFZxlZLb+hndZz
zFHI8iUhckXvLzwNXlX5TLC6TRZ8lsUj2IZN5abLptPLCfPCp7Wu+85UTj46
wixarl6a2K1JB61FiejFFrqtN9d0w6iDXnemg5yJFWZd/3eGpv+tpMjHdOnR
Ge3QGPlkEyS3QN2F+YyABhkHoUoXYxLPSEzWvQF5ChLe93nA4MKGwNqxBzuk
0D9lfMVKEMCNK9Ziffy0j86C+aiowMRaql23JkUS7eRXDxTgE6/4fDu9N0F7
jhD/3Unn1JM3zE/wdJ4ASKNkYdPOFMrrVtjdQT+A9Eakb95f9ExkEFb3QJTO
MrD84xTUFX5r3fkCCm2FvvHHNulR+PtAqyjTZYY73duC/+MPNzi7FWRaZ1ip
HnRk3SSmejzYrOLKh2HlLeOLJW5kw6A1eDnGhm221M4cOHSWF4sk3hxrypCi
1IXRR9Oq6IZqdI+JbkRjFazLpLIGkhfeG9CNk7iJjh5HBgmRURpCQdJIV2FC
WRqeU4g88HLtOTr8MRtBO8fqo5nCJ2V9X4YNfy5d/sFGsM8YNxBOp4UWJLKT
zzQX9nMMzvhkJFT4neZuDY4qmizX4pgL5hEBlHoAY/VQs86B8VPu6S0vSNb0
tFiRhSpXvMrJJZI3nqU//K/D5uul0IS5vzJL5QIVRCEj4m19yT8tliHI/iiz
z/hP+qAawPGHxRyONowRxlUSIVFo1L29wv9fEC0tkzAfW6ipSSMDBYYGMNOm
NZ2J5KnE70e0xU1r2tKpqLY9dzEHSHdBjqVkSrPh7Wn8u+oSGd8TWWgYLebs
B19k+M4+dZoY6sDRzXT0+lcniXmS3ZfanwrfbBzVkT6ViUE0izGfa8Dx+R6X
X2yLve6t+IsdUGn+7rgO49ornSoLijN9IBZDgllb2Jd0ccC8mm7EMRFLZH+V
22JgozO/X4OJdykbqljVv+NZ75AFQRPTwP4Y8UrF8eqi4efTTIxJ3i/pfB58
ByN4okL1BDLw8KcBz97A9SXK7e+tmhDrHFOVhiPc4Nd5HCIQRR2jghNaGDAI
SgEScCjnnzHLH93qv6noQ8idvrYF6djkztV7qKvQW+mf6AGnemRvQHjbl0r7
VfXGSvdGlY403HSwMfh+Lj6ulGu4yk1/21OcPcdLmTL0f31AuH/3MtsJBsZ4
D7tm4xVU8Y4NtnyDwAANxaP3Xng5Tv5arns6wvfiAbQ+0O3x6pfxBBdmuq0L
lGs41gZzQMI6RaL/jfDyA/E3++B3gxM5plThdVwspC/jisuln5nRpQXpCdHS
/nw+CMm2FEBVpV3n1p0987i7+ONLs/rcfqScFUiyg5zdZDSOE4GdRGT19XLY
WYT8fVnMyMccIaGgWXOzywQ3KlGd3MpG66bq54oVJBE3ObiFgrcA8dz/roLx
8WQR0AtRGQe+3mocaKJzChz9XSstq+v9xNWd5YJUK6HkEHzi52yNO58phzva
wPpMcJHnm6Hd5WojJpCPpubJW28s2w4tKTmR2Gkkrxp3ni21JYjGrYD1yffi
di2xfWFN+E0dUT1wN5q2iCXhd1f+CdCX9DGgagxrVVWh4yeVh6j4lWMnxOKk
r90WL/1/hQKh137a7c7K5m/UcfIuYxMQct2y5JCU94vdH/PaPg66uXhUho6s
pXMiBfLpdZxdeSD+u7RrjPbWaBuc+xIyv0YbLtcQaUyMDVoYNUjPoHXQKNGc
rw9cSzYIUGRTpFyDLsznzFDK1QE33P4ATePHreC4RkhMFZapU7qc0uRFmFZU
EoP01cfc5OxI6s2uhH97iT21go0fQaXxfvieBZj6bD9BC+rmdqonVn7EiIFa
yMAI23wMAwOzsdlIvlb6j61z4Z50Wrh7Jw9idUbHrImOaza4Xjg9VbkUq/Ya
OLLD+OumUKJNnYU5PnE9K3nsv13lIjqBZVYVlZD6O1tvO7HcqiFZrxcUl2k4
PVLNml+fJSMthCYSBtPtx8OLACTqVvNOBw9ALQT2Sx5EbZuZDRlJO4yBsD3B
7WJDLzZdHP6xNyEnMR63b7KSynd77cPy0MhpIkkfdLR+LzVidfSDWtobhQYw
htQbyWBMDHz5lZWKi542ZyvuJKaJI1z0Pb8SGX56Zpj5GxidS0EIvaeMOYdC
RD/6A4hSPVjuFsBOsOVr5nzpZOKkknH08liIc75wN2mxfUbZ7Kr4jeThpGag
XWmST/RuUxcodRO4KAh3IOFqwUrHG8L17d+OevG+g7Q8ypPpLx4fjjg5dOwf
hiQtxwNC1PDfAhBSeq/KXgaBSnEimYxJ6hZMLp/4YFzVMM9z7nwTR84B516d
H1hZ+PkwMw09OJNYgpKwBEla96jQNzyW0+h6Ypc8uavA8hkeryaqLgfm73eu
I6dymTqe1GlrmgSJWd0+pMvfT6nHaVTavln44kfYvfRJtTNZ1MeuhKAVM5ua
ndu1WDUrtRGcuPQ27np9HhLA0RigHYDws9NxzdtU/PozgPw02+QLZ3HWePzE
rspld/Stc8RudJvZnXslKB90X8/W5s+HfQq39sMtXNLUsssRZQVRASl7+5XH
pzGCdOGAcjCSdhf1Zf3SAsaC2aFfNUyqQNSZKBXhpibew1OaThu5AQAFuOnW
WOPIG3XCclL1SL5MnCCmfCe8jbP8iceJW/rghSIbsctzAGqR0eJtOJ2KMQBh
txWaY5C2uaSALti8CuLK9zSF3ql/zg7HXlYrZXnQ1HsTDcgy0iCT5MTqEmYG
9zOPxKQiF+a0zU0XZsy/SbWv5rklAWzTc4NQTqOBz7u935vLZkPeHJMQymsZ
YqQYzbdEGu7zpfl3XHbQep5X/XWGKi8GvOJJoMU2PQGt7jd0yrrXCMQejcUN
/GDRF7jCOWCo/Fc8Y5fT+asb6FWnuNOjAsHqo+2RzVkVfkxHE9NEM4jFWooS
Osfv2bnH2OVOI5wk7llUQ2MUyWjZXEtstLFAVshDE1jImz7ZC9JnbO7SbHlE
OEqgs0wtmOriUeqa2hZ8OF3xbIQ05EY/Tk3ENrardxpyptc8A8sWr8Xt37uT
MLTREiuiwnGuuuy7rtoFaAK5ogwxMiiREjKRGZuaKTTPNBKweUXpvgyeGM8p
8hauE0/mkpGv4fcZLaCeu/2BG+S2iNxzjMErQeFwsZIHCyXdDejRQm2lyM3g
BatzEswm+AUlqfbnYTtPgoMRGRskhQpI7RMAzlVvCFZQnWw5Ls3vcW7S2m80
w+auJ7e5i0KtBNxghsHuuY2mnIcva/qofHDUMtJHHbRx/s0j7fyb3HEiA4jH
ZMUe9mMmdBJGTLDYn+ujH/aeO+2AS4SyZ39dtBwx6cyDXc2RPOEpkMY1chsX
79IPIY0xM7+m43Tp9zVuNr0pZ9f7kOV0OoEO0INjW/cp0x+AGfuFnW4v/S+O
xo4ZtuoMLVBb3sKBZ8oIDcbH9ZMBAbMp40cngOVG+J7oMxe+BgzZ/kgNb1WG
1Q9k+HushilQzfBK9buXcqXP4M1JlpYcoRjsM+jv+pSLBXWTNLrq0FnpgENB
xYy16Wee3NQ8VabK30uNGMN8jC+kSjx4cQIcppqs9wT+Jf6sR7ZVShwlVxDK
zqhjTOQMSKuENrNHqDjr7nv8Crje2TVBo0PMaN+6MQ8xZY0ecx8XLe1BE8/P
ct/YfrjbkcAVtyO2pgpQtPnUHp6wJ+BIK5DU50hxVeZg2iO1QyHjMP1Hdggb
0OSkRz4X0hR2mwDX2dCdgYtLRY/KKf9JXV6xklM2OrJR0pHdPofQZjrVTJuc
0MwXN478ux1UXDLkC2yaMHha9VyAvjsKuz5Bq+oZTqf3eGX3tFLG6yS46hLT
91MY2TF2vz9VzujCXFrquzpj0mqDP7VwsUANYMyDbOV8n3dv5+qq1olPIqOg
REQlXYSi8waf+UbS8Jss8MN9X7u9YqYBhIuxeYa1VdF9sPJNc2CTJWsRLwTS
hqEegBOyjQQ+pgyxCFFFnYEr5MJPNellC6rFnVbT6Q3WhZB+eYmZ+pmSqLsz
TOYtluIlapQfjq9iKaax4gZIOodCFqyitvxBUaH1rEn/m4cC4VofcjNcuDjd
jXbBPzT0y7/15ToJ6dVod/XMLt0Hkox5FmflhnPngS5lWmuEyWn+MovU6QYz
wtJq+l765vpXtI9GUHqqQk+N+HIvN1KNZ8mXDrDrS/zIP815QD7Mi/yIYRoh
p7z6GwYFbPHlxVHYbjd9mZGAGVp4iGtAJ0WOE5gepQu1NJog8tiUKBhmgH4h
AKI2ul72/0pKtw4tqxix56adXHUH2uZ23AUXEaAych809Eg1RcJakgHaZ7+y
R0DT1Mu+lQXGN427NhnwmWK+vtugm+RGIGStMCDX/psDpwZmRkbubpLpJ0ky
6/QPJ1zubPK406Nki3LnCp7nqwKp4cogOWYAKTHvLOHRqH78fSiNZftJYoqf
jQVIjODgliviMcVg6BFJ4w0F/lohU4O7VCmpXc8PaKqMTNGm7S2M4zU6P2Dx
5A6CknyZyy8v1iMwF2tWjYmyFJmD7OcPR4g6AdX1jq1GBzJlo/RNH8gCHtD2
UJXEQKZ6R34Jwj2+s/jFOz5R/9sMsvdoBFee+zvoxFRvKWM5ttaMC3M1p/8s
pB1BChzCqUD42+dS8GxU3uPv42TnzuD5zYoOQFjdbfwyQqOI5dSl9xsjpcW5
yqDmPhNy0lInG8e8opEFQyrDFZI+KNE6NQWyMlaJAHgyfiKNPjL+d0iVKvGg
Mj47lFTRGKxc9gsbYEtJIGE21uNT7Dzl+fBxMpwGsNz6F56AgtFFTWvKzSW7
B7gSKBTE1ElsgwFhUvMAx2T0mahRLfWHuuimFkSmq53PEltI62GOodMgfLd/
Yh801JASHYs3Cd5IxoVXsElEVbC4vduTNrtcxq/PrXE95Nt+P2erDNhbt1Ur
MLNZ3lqlkqtHZRmkaHz0R5MNrYjQ651dX5OjYVtn1yTEYrXLUZe7cTu4WmfP
IT0PCUW4lLbAErTxyZMwkWB7khWkDKonjf2oA0oS9ampIDh/88azVYPKrcuw
kZw3TUMbGJGscnyJ9rVLh8MrErqxHJ6+URsx5ysf6xh5vkcJNqpl2xdi+324
8l8Z98nk71JVn9Ec0z5iXd8fHYZqdDC2S6Az9SawChc78M++ZuSbJ/G5ushC
pft7nyWRj/bcRW1TszZ2Izw8JkPg/nelHysmhDZeg+A7leOmWteihtJM8ktP
HCxRV4agFuiCwDavougkMR6YyJjVZsTRl7r3GQpI8/JQruXB9GQa93Aqq2Dc
o2VGinvzl46JA+yT8QKCIlmtkfl9dxktNjPZSrq/OlXpcl0ZZrB+ePiVOBRp
JeNWtHW0euWfSY5Q1mYOqgkUgZwFYuj82G5t02PUpx/xt6bEo/wZIaAkrHAi
HpchW/rVR5slZySBN606kRKKS9g+G1kioZfgpEHNWKQKYRTZUD7kljclSQwL
dPg6lzkdQlkIY/xZIw3442Zn/UFrWhwFXieCmi1sbqefLWIYg9MIRzurSLFZ
oYle5oWSCYcQ+YqsihlbHBKt/V5pXmZHI1i4UCO8Uhyz8K+7RsR+Mexcf4Ql
A3aLVKsQ4fInvFoGt+TwobFTPIHEcAbo0O62/Hvlu5eY9DUuXxW5Tmd8ZLp1
XSl5BOBHMEnU4DIcKZUmuxZ7/whqB/UUiNhpZVjGkN3T1vUH49IgYGp6gSB3
DtGmmtt+JtsF0/Lev230ytAFe3ReW7sC/fAX0gljPynsyuBVMJFiZY08C0E+
7/8MgmASgNb4y9atdIEkEIm/CbSjZK+zh2WO5j/R3DCCTExY3WFqhVXY5zxd
02Xli3AljqmjSdAqpONK773YrT8tuYT9BqwJalhRMjpqrdt5NO95jUy8znwK
8hDAbF/d6nsBCOKcWwomN1af6FqVSGvvFbnYXqD8ID6OzSmGqNG3Vzu9HQ1u
/h5yuR6GlHzGSXpusaXtLA1ZC+jRVf9lFJP5Ttn4yOR3TnXj7/7Z2k2I+UQZ
+ws0DjAcCPJAxYbiHm1njxhAWgl3JHrvCYNC6DLcot2mUUhxoaqm6yDi526K
WWiRMHM2qp/TCjJyJfvLzuvuFxgp1R0IFPb3DrOMWLUT/OXXIK1fXTL7BGuY
yMvpIQbD81DdsBpVoi1KOigHuHKFXc/8UTlc2sx/UBNaS4Jq65xZQJT7V5+m
5tmQ0HRw1TOL8rY0tXaKqPF4GVh+f8JlbDBL8fVv3ae4nlFE5aMZDWWVv6hz
fsJTl1m9bYYNOUblteTi7pkujm8pnrOwitoMvKuJPMLybV9SpaqUJIJiucnT
LDQv2rq3G9J4SOLjDDtHKMw0SGBanTz0YKvPJmXc7JWWokBFvxd5xSgwWB2A
DCzzQW4hpxEwdMTRPcLQBxGuxfCADnDSb0XCCjG0UpYXPP85/uWnTtCObzHS
e7L+W9idbkfpnZQuIr+j18augi1PG7LkjVlcxRHp4bEd9x8X/oEzjLBylXz7
7/LlWdBHXQdDG2v/AwMuApREM+Sh2ZV5MgfCOiF2yT4iuFZAvL1tYVjX7AAS
Mq4LHmj/wzSzbR8eGmEjToev6SbXZN5w8aWJ35RW1A0vCNN5gNdu5zWGDTl4
jFmFJzCJKv1YbRVRapxVraz4KXUkH2/Q0bWiVaymQjo4Z8E5AmIrWjG0VFU1
oYiZMhokt31Opi5n/HLnSWaS9o5ZKFOu1XIQtgf+OulIk1kXChGUbKBdKiFi
fwhzKM60bFQYzkm4BM+CEJFTg7MQ3vkE1rBKqCje39voY9CtlyC+Tz6+xcGy
ky18ZtGbXscVlosXHTwxlCNph+FprTxtfNbakF74py0OVPfMlj2UjdE4lXu+
sB6poKyrLbjHrR4NWvDZA6pRREkxuYGG5tTphJ5IrrCWQYBtI7evh9cA/8zi
HqYP7OEuXajMiHr//8g2nTCWRgwRyvxBFutO7WTCTm1NzApKGhKUh54wQd4U
R2re+sgJEhj2EFfKC/Y0OhFjvsWjjKHgZ002VIuYDhvbLt4VxpVngG8kcvOl
1vvqao6dAjG2hOFLHJxlvoLANQWlgNeP+LoNpPKkyITSoaExcINHREfJvb2/
Ug6AiqoQW/Kj2kdkuw+h7t9A1fwuzi8sNF+RryMjT8Kac0+nat001vez5S+g
ev88GxtlioWLb0kP9OaWSxVrkD+deFj/ADgkWqoX/FmTG1HbgdsAgbtph4rZ
25Yn+ErQpsww1Na/d7aVXaU64DfyxNs5+UIHyCX+NWmRyYOMsYgOEZgTCuli
jraJdHBlGAp72kl4iOsbybbRylxcjH2mmwo0DuEqPwGrV9upVmoi2pFl7+xa
a/Uce3w21F8iSdu3/QAu88Btw0t7efacqdOLN9bTh8aKWCAZuV3ju1ZqAzCt
ho1VOj6q5heo81Kq6UnSLMgIZ7pFm1iCiJaSB+uiHe59cUly7n/qi545dRmz
Y8e4C9rjcabBqWyd/5hRh2+e8TpdLEkh4cEOInIG80+J929vw7ChlWPITc2t
32Vu1MSSfUQRQu7kMC+NjD4WDvrFFYqFb4NS0CgHFY10Fz3zrQLXAdfwKRVp
iRDXII2Kb6Q0xdEubvXR5IY9cmeg6iFh25CXJrOi/UG62T8jKCHpl/MBisqK
eE8S+4QEVpsVr2MLmAvlRRXOGBg4BnER1w3J3Y6FbO+tdvK47xTYe92rL8bg
qGBumuxGcikenmDco+8FhkrSV0W233Lq2Qbk1HbirHuv8EKX93DdY+YKtcHC
pPi4RJ/7hBmESvu+G2Wpor4v/T8xZxzVTIpNkP4mia11sSQbDc1h8iZoHtdB
8Q1VizfLrIpGPNdJRdNiXy8ErvPmn37VL+Zx/RoAAA+G1TElnhZIfJOMmD5R
vKoHpkuX26U4FYKtdhURilZd47hy9HkoQlHk8mGFj+mdY78EwCNr6vmBXW33
06tvhEA7JfMXDzMNdz1AXMLbe9tGbaOL5vyfjyJYSxwY3ffseqhYWkqCo4OF
qDbwb0ZmfeZ38qr6VA/APgnrwGPl3HHJjVczzPsxx99F+8uOTT8JGANMpK41
W1AsNZ88NRaqa4Yz2r8y2nULdPYtPcqlmxjdymsLvm1M+hXhcmiTkFcZ5aeD
1JCS30BSwUDx+4DMSFnajidguMRlqEd0B5wEWdwvqiLuiyngNkEEV8Ak9nMX
Hq3++VmLZwDRT8cBdbIEQgPf+rTy5ffkUqi7Q830Daz0pYGn13ZMRm/QEPmS
jKw9ehuq9g9wbooiRvTkiUYSmZPc88clx1JynH9jITYZaluyFD2saCfSUQfo
8+vyb+HQQ9AaxQMRsJiZ8kQxRCel85fDYiO4oX+3u8oz427eE1Cfs6XRlNi3
fbKT5qGTufoT1rDWzGQOgdNXOngRy2Q2FCxxwsFUOnq/wAw0yeOwOgPycjRj
rDcsPlPNfiCph66Tx6mucZgMHKEn4U/Os/NBGWljzqoLBpZhlXR5TLfQDSnk
1aLLV/x3sBA0CM5IvU9XCCKyqmkTYY3Ay+jBCFYD+tWtnKDjTQ6EUcogoT8L
EkDqZHKYrea6W2MZYvNQOHMAtPXImBAsoE1tr4jC64NmWyenVjBTtTZYGGpw
/uIfQ5GoYd1EJrdbVlrpjTw2JlAlYPUWqNN9cayGgY/XBRuIvYRoWGguuRny
zyKbwt7rfiEjDDZAMWHoADEOwxIacwGPSfXcpYwL0rAlsLge8ecP4S5HSxvN
FXYdpPtXq0FSe9X7GmoEtoZKo6OqwVB2YF/ulYj8wv2pIokmn93Hcc4ZCGRq
VoRKavWLj3cNXzEsKKLu6kJAMqz1geWUQ5mImc/9E7P0XZs2P2d1aK/jinaM
q5Wf7T1i6WKv4/K76GWEMplKLh0CvAJTg9I7T6q+rNplWv2ade0QV7ne6h3h
WIwJSyJPUzGbc0ZiwZ4rr/McodblYe5CEXs6nGF8uf61nDov44M9CVk64Iux
BxGI2Kd/oFmycEVH/j61+KeRXR6u5qoChewxGpzVK3LfvhPutp/17mbLKxjg
eV4mktLpWNflpevRmpG3X9R4TNoUx4AwUmHGLtvqFbvy5FNXhTJfmMvTTD/t
iJeHuu7/mXdLG0stiqmqGYsRKVTVecEjwG6j3dimYBtipNc+Ft/JJAk03i3I
0x3D0lS9us2j5SXVO3qWECn0SqCtaeK9qUDe9699BTqhp6/MRz8B6AXiZ3SO
JYQpsnWVtk9WCPJ0QEPr7XEkyV+SMgFmrP169GgQaL/GQV7+e5ZywweNc4k+
75kt5grOo6CfPoJ/tIm7U/RvFJCLRpcsWIyyJUZeLGmRZrt1cwEu+3LHm7aX
vbEfV215UR9tP3dHS95XARvWR41hVu2jWHn+XCahnMgA571ctGFUHB4PUkTo
kInaWVq0cbsDUkt2jkY9Jrfgdpts8+s8OVoRh/ZApFwrcYj6ZV0SjKdbEY/P
Ndh63ixcxyKP0k5KZnz0Q8WehBCanVX3FyJaM2n7dAC3y8vBpCmtT5t/zmmC
JQZtdw9/eXHIrkY7j91cchEItCfXou+zu30jqFHeW5jNVE+R+OrtgSO84ifC
TWbTEYi5OEtWB6RT3C0v5v/i49I9vpoCTI4YLtn4xqFRj5T/etWHZb76z6su
lAJNDNYJuo3v5lP5QalI7MFAutfWkg/RTBomvWQEh826qwKwFYko1udscuFx
GYuN3SovCdwfclmo1B4N+A8qH7Dq64euiAKjPkpsjvfL02Q4A5mAKezgUCmI
/Q5iT/nL0DFcoH8fVDMbLG+eutNP1s/N1jnu94g5LBUR9mh+6cFdj/ChbvIn
FyON5LPeSNunACNieMprnqEMhi0OGfe5jsghQpj3mR9tGTbN6Pa7PCpHLION
OQcwIY4vVUhq8KuBV+uA0MZR6sGrUcN0usMAL/fwwkw/R1AX4tqX/Si2e8et
k3QzWx0HrXjgpkBnOCCYPm5R7encv9vJHUtcbd7l5nV3SArHjg/bM4hgxRH6
dvGT9yarP3dPSD8fShJwImEUfHOob2FtBe2oiFoCvsKtkQuZDfHNdo3T4Eaq
m3kIXKcJX718Bolv+d0VLOUqH3eWQA7kUXUbOYkSsExOVa890DBA1MT45A90
Xq9SPPhky9nECQ3MAnzGzgHwb5ZhDZXDZu3qKEKoq5Whf71/SrTeRiDXg/ey
uS60zy2MgMsltkiz4lVslZ/LuPXlM3hOQ2v1380VAzEG6XNTBqoET+D6jrjo
CSKDe3h7biQNUUaiTsu1RNoSP6OUXFM/ykXNZcB4uta73chLFbxqw3X6CxGd
cmO5PuFedvvfKxvb/rx3/tGW5IYVtchOlChyBVSZbPiPPPqs9pQ5g3hUCnMg
DvY37wPAc0J/TJ2+04tVaDWRlQXDoS+JcVg7nm+lcCEmbRfoLtXqz2yusQla
LDiW352GOKpJ9LSjgaUjNPghA+sqiCbtAIajdJiblhqa6qH4XmKplkNPkOTd
vBF+Wrh/99/gdjSj3NCIa16EWxZdiQpwBaUrMRlPY8ZtmMloGxNUNVIkj7ML
bE2MoNf0PrjRqXqEyNm2UZjHt45U/vrWRfbzC7f124T6ULg+gGDIx0R+fhPC
gUWoC4SbmZZTmR4uUB1MiMopmf3pezXNfloYWdMpsgufjGqQyrmKwr8ugtZC
Z5eGb3rjcWWPFZiEzVWIFsOh8y1is3kkCxCCbmmp60UsJ55uLMNcXjM2SsPJ
YzNXOAPUnOzOI9ULkoI7OecGzre0s9htRa0e/+cJ9ux6jYYYPWunpazCK9B8
rdL4SfyGP1/arlhAGcNzEWrFMlH5D/JKh6lIijc0lx7UEB9COM7tBLiY/hfY
xtHDEnoBHMGXc6usKrEt+utxXpobD2Vfz64ilvagv6V+FsTmCGRC3tn0/wHG
VDgFjgLMXvp+0nwvaOfWH8MGuQQi1Ksi3XyKCZ8tacLRbNYuDx0an6kLREv+
6CtcHdiaM5GXcHBjBStC+QgJkEhVzdB47Qr/9qz0Aeb4iEwwP4rBHQSA4oXY
wO2P9/IPoOe9MVeMH/qECMxOaTl7RnJGDMH0bUhtmMtCisj2J3s7NC9ojnA0
tTKeArA/dOg3tJFe0wwYZtH7CVfFdWoC2clUjYSieyRbD5FcDy4ZGr9tTGDH
hv8TPN77/1q8SwmbH0OZM8yK2s7jlRlJsQtkltK5iWgHXoCwadKVFQacuRfB
+5y3X4HJkDp2PHsfpG4TAnSYvFYx66xfQy9LuJobjHq41uhc5NdWsyPfwRzW
OvoMGwqWYlLOWGLy2t+bJ/IQO9riqxWCJ08ozLNN68Kw6qGqfJqcPww3Pevk
BygdbEyvG17yUU7pi07FVKxbbuoYve9xgHyHVCFule3pxNSKIADd63B2HSr4
YjBqSQX1mCpwFITEWn6/uK2r0CPMzYxD+XaomrgjEkO7vU0LpuAgXryx9Kde
BHoNzBMtBOFNGmANbX9wFwCaZ9/xQG9CobtckW+z/m70aWW5i5LYSyzsq/qs
hOuSfZJ0Sq+6gULvSX2TP8Rk12Kp3UUhFg2lqJ2TlV/aNuOCDlr6Q3rwHm0u
yPoWwiM7/jk+Xs13c2OVWq+9i6viLZpHKiOlxiK6aXoWG3ZtHJk+ga04q1/j
PsU3QUlHsFeQ+I4Df5PeLTewfxYFF85aiQqw7Fa43Mz4+ANwQ8QHH8pPlPjw
pqv99zH1fQabngQpKNjKhdQP0hKxZ+CG5LDiXXDAsBi0ITQ8eNVFZZ07V0p8
w4FZ2uNfl38TIdhH0TIxicpNmd0C4oQ+VZppGq7NZxUABC/vix2frZFEnALH
v29um3rpFDG8B6Fb7INKENBg2xWV4o1QDI16dsk3/UACT7coyxRd5zKO5VVo
Bwss/PLMWpEuU067l8Ow+uSFSiShrbDsDRdFOvoULF2iLrb5AisGWtYwgxvP
OQFU37d2CynvhB5IUoeYppOlL3Tc8OM3VSGWCmRSRwDwkctmHsJJflULFqtl
32+6IbeWCR8j5DhnARbbUitD2sF8tfNCfgZjSBbhj9SAsu0h9rxyHsy9o5WQ
3uLZmK49Cfsr3qa7XKHGMK6LnDIEmYVUikqYmoHzF71jHf7AepM8ccFQMO4J
MDb01P7p13SJaCkDQU4v8jjtwsk1qIskT/svwccBogsFySNQUaEAxtmfZc/y
TLL/0FW0UW7K6cjr3Q5ubt3qmzdpjS+TLdjW77cq4/3EPMRbMCJLka/9DdJR
jDhIhU6YuXsvhGf1hSItIPMJkgReVdOQIpe8DpGdousixnn/xpEZkjjMgFEZ
NSZ+sfWvqndXJLXbGJ1jS50QfgWxwCmRIcRlpkom6y2PEC7lAZ2GIph4mLRW
zTlqEN/j+wPGYBKIjDc1z5K+WdH20+0DYmH+iEdNyj95Hiw9WOhZVwVDxLNP
X3gIx3nvoiHH4PvoKSAR0kvT6ujQuxUpwhWoHdD+v75j0v7f7nJAMKSaJmNG
4p9fQ6M44kinfEFsmr8oIEkHmLQ0+QVRNDId/OT/S1MxhkHNd9hSIEg0rYcv
H2ul7KY1MDZlSyzedF16ghrB5VgfPUVr/dZZV4ltAX1wGS8UVLnneT/uYHZI
XRFJqt0GLyLMV4UwuSY9TNe7M0aqLNMYqK1wUz2wXAn9YNAYwcvOXqPhu7hd
D0R+M5TGxoyopVJ1WjO8lmU08CjOXDzeo/3j0mn1ZL0J80+GOpl41J5Vgp6v
3hmBwFsWlcbPYicIJrRx5jq+X5bzhDgATbuHdkndHZAIf4D11nz1ZtrJYXVH
ffD/MTByig2aQy8l9ukZR+x5G7OKXdglp3thDS9Tqp/idOEY24yeNqHXtnwP
lsq+GgbvJxBp02KHiE4YwmkjvFh2vSjxzXT8YfmtiBXlWhg1eJTD498gizwA
XZgMGSEg3F/au6XxWvLnlN/wDYIYvBASIfyZiPdbWlVaReZDtHCVEaVE6CDT
K4bcZFVql3d7Yr3KY71UME+2VV9ArJAUtfj6cCU2kkOpg/iAiRjPFnTjTYTv
n8pQjf/Pb9oeHnlh/v/+mDgXzvMHvdPFHNyPRot33T12ZrOARotodtCsthJS
hK6GW4KukMV0yHF+BY0KoSqwewfHFoi0f1fSjXns9BcJV1IBgnXIFvjR8KoL
EOkQ+ess9YWSZekbC7BsO5Hj+XluR/K1+rabdsMbfbrSSwT1WciJLfwwRjH+
8PPxQMjAZsfrD5mcLnzNcpKhmT63HV2PU4Svkrr/6m3VmG0145AY7JMgxF1G
nsZMd9lzGGkoV/pJRJiB2BAJn7yHiZ46EnzLXRCzzeds1c5d1BHd+ejkJIk8
DQ06UzZFrPMOj9CV+QyCiMYVrwjRW7bxqdTZ4VL6X7C0XaHaYlrbl3giKP3m
5ipMzpiVmuOwB4pIc2tkp4lDcAw5reHY2zriVkO05Cxj0lands0Kg41s8W5O
c6xZWkj4m1Vyi/ZDn4lIp/3BxbuRzAVkdVj/jcjtR6l07m/8sFOcMVnC1kK8
Jc3XPcAWBvbWo2TiHplTF0QcZVJNgc9trGJkuk9vU/WG+Cb2eIat9H+iZx4N
Hu/zIpN/yrjslIKfM/MHwHdgXqucuclbE6DKh0Zx0ly9/pgKcOKcRTUDRaec
6qrNx9tC9kEvNBS33pVqM7Tzf1BQYS82rdePJ2tXmMctVo0dlU5SvpHmJwK/
SeFA47RL14Vd1smXwdjeaOMUli0xnVx8nNZVj3/JUDBLMQKdSLIVjIuJl090
npDJpmv0It1VUhTx5MT+YEVr3/IlstQX2Kq3oubfh21aImtN1wK3bs6dmPm+
PfjjPhrhLaBeb69wdLdpx6CHJ6OhwzOBH8agDRJbqqGd4bc2YkgP5xZNLJdI
EcVp67Gc0AYtE6NZuklnYH/OlXlYa+jb18sUTPN5H++1PDDHIRRKdW6hcQv1
ID2ZeOdPWxnmWfLNtdcOX9I4wGrKm63QS4QKtQjJELXodcErAlzP42iKZuJX
WLZ6TMobDk2uG+10Rt5v1RLKDc1i1SYx9k0nsgXkj9slYAK2AFi1XqcmKwqQ
LtQ8UJtr66OsEyDikui/xe3V+alVB25z1bB8r0yF3VXQPVW2hskZlE/xr6Te
mg3vdjmn+6XmvfxlTSRY64D7GC3iBF0Rm/9rQ5Jkfczz7gJBlU4maxk3T1/n
K58eb/q777MQtfgqkazox9qC7z/buqj43AFySXJ5eOaN0e1iPS16xEyl2qu4
aEGboiBeG+0TAd0ZkOSVSGnohRPdIsxN+EaMZq5v4RLeT72VXxGwLjEo/AVu
SgAqK19ohLACr8++nJ3YrE3ZUus6u7JIjyPox5+K3tZgjQqCV02mjRplu/Bu
qXrPBCpz3NfTFVq7YPs/0wJP/nHJu7L5kV2eCuzN2vDtfkuZQzV25SlIps7x
fFkfM/47ZpLwb7UlBSWPLxA711Bo2XpQJsPw+5qbIKUL+jvUAzsj3Eay6mhm
xFSrh2cZBMKF3dHyGu+/y5UA77DgMnvgeiFEsN85WwoHp3WuxMHrJdrU4dal
nMv+zRbBr9HGncsBH6yq59g2232HxP+Db74ZP2C0cKqIJ2YnK3CQhOhRUlJ2
9DbTMxfHUMHgK0Tmq9mcpMW98FEV04nq5HRFINmLxFU0Zl0sd4B4E+7guMJr
xBFuLlQ+/dkWuMmCCgAvNFkSrVLs6l0gbrzQecy/as+IZXBFl8Thl5+QCsOY
dzkelnBQJjqwK94Ojo23bewa19kLwbTKW2gJ4140YXaO8eqXDc1MRyARmnq1
/I0pLFd2F2bExsBIpe90Dp1F6oYivSEZKdZfnqqzaH82OGrarzYPkWzqff2w
to6o98URWNm/MK8/Px4iIFulx2kfWRn4jE6YM1GybLL9BpCbe1FOpQaPjZk0
5RyN61LEQTGfdXV3DYDBfLa1dQati2UxeBYC5DEauixXR90hrQ+vX2cQ4scB
bRynaEs0/rMba6pjIhxZO7lkEmTvh79Qv3yAeCojSKUB+xYh8ysopfI16SJC
EsxnC2TaEmZJDsiqwzrFKRe5C8BZibJaGBDrFd9yox8dbrxKeMYjPSAeNynR
UO39+UD8cMJCrRHMVqiL+OAMGJdUA1bh7YBPxMim5qD2OtYmTCWS+iFJYJYx
JitcYLUM0tZ4iZWv4VCzrdJFyjD/uGidUox31AYCTzT3qEwF2Y3YT8FBek9O
0GDcMbld0O1X/6zZ+E3dIwG5nkBIMltA5sYcN3/71DR3YG0ExZ/kmSK8W1F8
ctxB71/lCWv/COcTWVSMPGIMgNxqJ6iPkWAypRn++nrrCARAJj/5cMfP+Nzu
MCex7Ie3OlT8Kk0DCtH6r3ZbZIa2QczS3tRKBKmGtxtFIP1FKMvZDHYxI++0
WjN8dcsTrSEr5e5EVGgP+oxm5lRV8iMkVcOlYRN55VQpA9Byv25Jtw6piKrJ
IN/FUUyVkTuyQ5NZDT+hf+zo5S/dxmPTvmcqNVnUUTCloT+WE36hFUA70e7h
LXG+xpwcuOfQzhzMnPKG8eH/kRpsmkej31iDN2s8JvtMbia2rnD7TwN4emRk
NwP5pN2gf/bnsR31JjUP6q0AhdsBo6Daml9L/Pc8IZ+FIGxILhZjMMnn83Sy
trB4hHW5hUkdhnfJ9mzncOBHr1cDjhooLEC+yE0xas0BvzAnwelDqGWAbonk
AvBqoFa3aKocv9Ucu7LzEkbMqqz0/7F9YBT2QPq7v0lSoYdY9MoY2vWmM3BX
mzp9xGkAxKGZDUI663HSSPuiYhhpHuxCWBMr8yDtzuhITmT+Sar5rw0x+bxg
qUsqDhpDAyCFRSk385Zwn7uKZ9O/dtAdfVJBxfHHVMLeIzl8ekFRxjwdOJm9
Ilh4KpHIT8PkkiBtkM5LPKBwBMYiFgSC/iN17mgN5uL/bmPDETRPCaOixUVJ
1njwkRozrIC1IumBRnjqwwibaQSvSuXJhh/PpD4Mq3klYZyDvKf3q9w1WJRN
6h7ot5RRMuJ/Dy47CW/GAllZWc2PsH8FljK57KWEqgObOOMuVPTwrbTVpOpF
suYigDWdHGmRCprAzAmLpu2IRF0Gm8QObClUs9ATxqqex6aXbIEktO+k5C6t
6Y17jIfuFddsNJoyoIAAlKlJWO1ETHWyAX5h//RMH8QEiorb9uJwl7a99ZCq
3uPwV0l2fwgYhZ4gEvDStoaEzHzuM2/r/UjqiZ46AeH611coRVZ97ufp9X2S
Apxrsn7VotfNTANFfNN87oXbZ0guKuynef9eDqUIYyOKDUJKnc1/yT0uhzZi
HDVGs0X+DYTx55vpknC0dybLpKpkfkCTA+T7LkG3PkuTk8n610aEI/jxx9pG
EDFz37q1bOwxdgDao0JbCQAIHdECpQ05sZi4iLvUOKwiTu/da3AVTo45ppXU
OQw7BZSN1N9dJT6lYAWbuGujDEgEsrJcsVnZGwkW5ZIpQ0GNiXK4sL9D00Q1
qKS9JkMXxzsj014jxSyUEJ+xQk+uAqWP+wEzhBB53T3oGHscmGWtro+D2o7j
xr8rtPo69SiDdb5DVxVisWo77nLVhOLKyVyPMG9Jex5ckijsQ46MJGfs8VsK
y6PYBV+BuSo8zCoUhYxyfB5XCVBD4zP91xcWJ/KNJ5N7tOm7jZK22hyIOdeC
3MEtdJY6jaD2rWm4aQouB56buuAI04r2nhuYg6Lq5Di7A3oKz5ck+IKijHam
xdZ5mKA1Jgr9noPdKXv9XBacrMx1f2hsmv9EWKig87ViA4nz0FJWzQo273Q6
cZeOg9aQM8SqEq8NAv79Vcn+IUbYLCQ97LFmNEKKL5PMkcm9vrlJrlv359EC
OKmUi8clnIjuGRkwIYsq3zAi0JuPHuR9isR0M4nse/3zXKe+zjpZMLmaMALF
id5gGj3/qCmXO2EmuW7W9dNAMvCvcg4izhBflBfhByKOqsRV/iR28L6zgg2e
IQPgFYw/OAQ8Fup26jgZ7OduTfmTaJVBOP8Q7tEUCDe8UY9l4oYdxM/Ns37R
HSOchKl18x8aG9QCRTIXWLvj1+tMiVeJ3+ObF/jDvwgVxGILjMNu8I+pNKb/
HTvh+FNc392eD7cHZtFJE0s0FInBQ7sroBdIWGs2/pcNtxPbkt/CZJaaUDpr
j0bhdDnwlUYWLTcw7q/lx7OfZeljkfKQd+HJ1smd0XgdzP02qmiq1Yl09znQ
sGe3wzpyXhi/srb/fsgmhohtKwQZj0mEkwgTEKuxUvdX582EvP3KBPCURUw6
eVlW+tYfLUqR9bcxOq31Z0jO6eLOuU9ASNL1lV4WTamVs4Bogrn1atRe9URX
2GhR7/yFhjMuuNvuthzXS9IRiE7/mjAp9eEhQfjJkZNE9xyHEA5vA8/DV4us
xsu2pu+IvlIW68ZBmmRBjshhL8UnTkb2oey7wZiEfDQ8w4Q108vYRuUd7Z1g
d66IQQ4vlYUBBQQT1PFrPl3d6bYeHG0vPhMeHemp3c/cPbFrTGI9hkwdn3BQ
MTg8s53rGKWhbbsAfguN8G3t8TiGg8KN2BfAoNncc5Wbc514FPHTxPX9LVXc
nyinA2HFIEhWg8VbjPkRs5WZCtTtuv1ISQSmdLHTOuVc/VH4D9z2tAaEJylN
l0p5t4bVIZoBG+/cqloIMVgSmfTvGexwTGOfgyyzcL2KSC1hlT15h948FyZP
VIojxUpKCVBEJ8sdbVFgOHtVqYVp2BXcaCmaYZAdARL8G5aIEIo3PPDceDJo
cEAwRqFTVTAXqDLNEAva0Uu7kEpDXtMCFdqJuTpMii/i1lafOa7ot+aToVd8
onW5jtLvbL3sxPko9SwjSsEscVEnZazt1BVneGKyCkDIIa11pMVoi/trNrw6
Q/hq2kvUv8eMyBSrP2117A2ZMEuW88BiY2dCpIF3HK8g/Wi3Oa+GVdn14/e0
Evw2u5f/RWtLXo1EG6kwPSwRVvV7AkDer73IK1mM2euddrJo+ieckig1Gqj7
/XOl5Oik5hCX9pLUWRdNu3iDZuHF2ORWCSO4BRiH9bq+96ON1D+SzcNNeCm3
ctYDx7y6alxkyghsDdtW57pvZ3vEDMqNuoOl/gxqj5PltpYKUJj4RdNMDGPw
7qJTYU+zYV3oV0ZouJPaXOc8+0D1CHaXsRhzqk6nKW6IPL2/Tbl7dmYf0GEK
xdfrF7K1h4SF+bv23D2JN4QxwBhOfj+LydSsruuqULU4p65TgrPpMOd0zalF
gaw7lKh1JogkUAtx4xUhNoHLUDPfJbeDCFOr8U9fS4kXDK2NetikxZ7IkSRc
H796OK8asOKRzebItwNd9OHqC+cIU6GF29kC1qkpR49qQE6eNefCGdEiEy/7
M6Ti+M/Tq9SW4ww3VuJD+cU9wTcN1pxahrkG16/7JSrQeniusSF73pMXp3cq
sSRL1+mWo/QjgIpxbtbmPIl3UdVcHYUNn+rjMuD7klnoh5+E3eUh3Os6FSQd
LCFxZx1yHuqXAFcAUybQdHNpQfwCzPmScRywficPltZh5OClIPbULqQ4FcpY
U4PiBlMMdRgQSxWpDAPfnKltoWnjqihgrIl9Q4rpoM6vN8TuyolJa1eIjBao
XcVuNukHU6R13OGQ8ZC3AzSCPtKTt1AqdlaGLRsmA/nQA88M4JAFvMVq+naZ
whvD/vVqlYXW1WPmWN7QOZGGM07oJ4rmXqgahmFsz5xngHSs6tw05jKMwC74
z7L6ZE6V0OAxo5ahKoXc73nxg7jfAfw9VaR3iUeY3VYlyEwe6N+zlg6WV3UM
cIFp37E3AqiOKEsE/Za3k7ULQYewmkyLtPm2lZDVBRYw8xaLzgOK1bvmCC3M
hz/Hx/vhP3PbMVgShFlPbtiDy9dAmkK8VGEVo9LKUdPlLEbJV5MBPs8F4nJx
Q/uKxu7+AymHy7UgsEbVaiy5gZDYabaVKjzoDRRb5QdT2MxMMd/O4Ll9HNsP
BbHHo3ND7XVIQHTT+mhF7wdEqKlvNracmIY1nuJxLTLhjs5qomo8svGujp1d
nZIOIQ+DBz7o8xxOyGqgvbemzJKKW/AFTFCNealXAc1wRpR6RF8v1wHdli54
LCU5Fg/1voW9rnNuYBar9XJwFcw5hhgaTHvH7X3Q4dC+nKszkbkXlHlnxxDb
3Nx2Y8L2YbNkrI8ljE1Ox14n7A0qa5trV4qTgbACx6x3gaxsjPjirBnEwps9
7Vkk7rKJWBHgpqAsSNEIwvdpLsdUIJrbPBmfVhI2UE6ZgZRtsp4f7f29V7HG
inbEuzcu9sK7F6+BM2tpmmQu2sgZ0E4MIrNzz5ho4nVPy+QBXLHOmjkXydEn
MWPU522ZJ0kAYsno2jd0Yf7+NLeB9JXW7T5YVdX5OL8AektlFsTV16d6FUPJ
KxhRWjpk5X+dxp/0VGSToGCAqJMO04V4QEnb9Yv6oZssopPoCfJSFuWe/iTw
M0Kyc91vgJXd1Jgqj+8UD5FJYVaurCcbdZcDWxBV07ZjEPwmsH/EyDcDIlmp
umCLSD2c7/xZUBZk9+INkDfFsPDJf4Uh9OuccHGRQIfTOTFC2G5ZtznVzsZo
E+vWHBlJzQGFXyCOTSTK7BgHubT0j/Y/n7HZC54x9PZxL0eRp5X4RzruEAGw
Ep9Ea6upZQIlZnFHYQYo2zSOm0fLTNkwceKnGxVdH7qXo/iZyuYZVjM05RGi
Xs+9HN6xGUXa2Z8TzTLqiIRuSnjqEcA/gCAT3H/5nV3t1v8j/TtZ+D5tFovj
CEp+Gm8hr0dbBDzoLpWZQX0PNsHHDoWYkIOCfRLPcL1QcVyMwUqi116TtTaa
TVj0DffE8rU9BOZMH4md8eKmx+OQs2eNlTchzrQKWjFMz/+ZHCQlBH3AWbu6
zehCJ4mhJ1JU6qLbnILzpi00sJV8tj/nOYxY9+yAumG0s2r0HWxntpu0dwOh
3TLpvwCXVKbBuirEVi04IA0jA8FwLNrP1XX7qs6tK8/NpBqTc8maGdnx4UvL
ZIQzyc1ucKHVqxMH17MVpIgJ5wXCDYviKAJ2OqKEoIzCSLYN7cNstmY4lcVJ
Oz93semxuKk3OPP6i3+AGK5XrTmd2yX9AQM0OrwuZa0z+ah49bl6rqr/Mvjc
Q/WOO4PFjgDz21hApyLpAQZvgfEsRaBdpwDClQsGYFTYuOoP2V5EU1beCNao
+mK31/wyevn3LRNVeiX8RQry1m3y+Y2WxTtyzW8WDwKxk7PW19yA87Gem4lA
tz93khWU2ZIDvpZnG3q/Gd8cl9lzoBASEt9XpufrfjVRzpH3Q/JfMAQLyPWr
16ErcSztOcJ+CTcB9GAu5NIqSRUK9GNezhquwQUP634JqZ8NxSdUXWNB970u
VBiQDVO4ik5kSxfM0rbdDTSGjUQVM9nBtHXzzmmckiZxMmtRPh9Sd2n51Hbu
r2iBHa5hAveLWzGm2ptLTGunE69NRf6UyH+Zxgef3l6wzBykpNVh4zL4NwKO
fUvrkJelmrchHzAjc7r7K/Cj+mOFimRyAM1h6ub9Qs+8t7LmF5ORsErX5kiT
u8OVdio2Zp8IVl2SoyxTipwAMnGaZSfl+oeH9KVdDem+n51k4ytGnid5doyX
ucUe5XBB26AmMCxx0Iouqj/2XKQGWjiSuuIfEMv4pEpRzujAiacuUIuIoIaF
D5BclLIOecBAk16izrEohmV9xoNO9XB3Eh2LY1cGqGWel2vb06mXYcpXKKRk
hvzZzfYrjznxFVPq9npmlpkOwrUq3LQu9cG3W3DxgNLuqt8uVervvlefyKVG
1BrJeZr35ZkFO7z6xNvzZDpIpHbITBvmu0le6VSAq2bwfuRjqmkXd3DsCIwL
+3PPj8NRtQoge8XwPwghoNmZLnY9PvoZqh6XYqQ4hLCJAmPV/nTGdfS0j3V6
wZfwOf1PNUSdS9rd4o3Agc5741B6OkdpykGFXp6TJYBx/L+XYtkceaf7/hBq
zZUOJaV0F4rxXCg8DPTcvKB0F3eLKTPOfmpwcnWjCQtoS4d7PGvB0rRH5bTq
Lo26b72l0z8//0WjcjjJoqKcrzVJ5nU0LaM/buk8NJ7JSpLKtADDg5epTVVL
A4yZzGXTcJ7wcTt3DxpFCAld2F2K6X0qV9tmw8ivNPzjMk96rSZiwCo6m+AT
+WxCq82VUAKxuwV6/aqodQql0OcS8EaiuGJL+9oPJYrPC+AMA8za99pne0S3
LZexkF7vloON5cuIkHV6h6CsBHPfmLnKWYkmI6fi+4M7iJii4UibWOG+Aox6
MkE8pFof9tq6NYtmwa2cmewQp+vxUJhtEYb5vVpBKd/fPRP4I90mhoEc6N1f
zICbws5GJRur/fN6/fb1bTtyKrlxpNjNstXtx82TsB6+ZdfLdE9BlhGJzcJk
Ei3sgQsTALlkWDPYucuVe9ZD3agTbP7RsFSNgvuOtDt4NfQGtgX61RKJFhEs
b5tJ76uRJwGT3zpeBftzc6zjbIaLJgHbPVXRUtkRA/h4zFyJ7MXx22mxb3Q7
myat4fgU5FSiN/QYQybHDtpEgE4uRDaWXYNmijHZOj9VXLn8zv63t6xGWnYZ
5TXbLmUeFBZAWQDaft4H8sP9s6BNT+ipAriguluyX9yhR8T14Vq30E+38Mpr
GmehGDerNtT8yaYR4USzVOOdXNTmBq55igtp84D8VZWUuUlqmMT22hGh7opp
Y+40kOuHiqXlDMVRVY32qxzxe13OcTh2WvniyIvD6UFx3unDUYt5D/odzVeJ
9heyjiDO2gUI26z1bglZDPCE+q6zPrxHhTpeXsWqRLG/tH/7VBhnHxKjvX7+
PCqBSqlEhaMTyAwr9c1b0ZhBkXddo6pD/+EEPQ95GX3Y7Cr2f/DYFTRILpUC
KIPMCVKxGYlApY3v5Y3I2YZy1NVlNvtkQ08wnk0tvs0u/GkLqGCO121wC17m
4SgyK/2wobDL6J1NvzUr7b1HzUJAxAjMY/0i451VA80C88Y6XibAj3u2LxZ/
fT4ivfnYPL20VKXC6Oww3xRoB7Ih9f6T44jQIUTl4ni/C3IWjFz9RhNvep3g
FDRHjffLy46uv8GYlh+8g5UkCeVtTd2c7GUARhhc9UshDdOf8mzzZ4BWm2/e
8dwzLEV0UEh/H7LxwHs3/h2pAJ3N8wXOiTATf2TiCFPHsaiF/YT7ZCg8W9d/
jHIAjr6+4v1uvkt7Hv9YEvUi+ieAHrA7oEeB1sTErOk2XdTC0nJIiYyKFCYC
DEy6lxAIQeT1xwchsvGRjjs8RVP3HXGz4aqTIEmu/L3XzoFYT5AO5VI6ZZhr
wfMUYfAu5ybjVWw8u1vrl6p3Isc/F2nf0TSFOyu4sNIyUb846W4EX961VGIX
Sj+adVfIxSgMIVXET6e+ZifMeKJP9xQKSGItmI8kIhw4/gx933iQ3TfSEOCL
JqG31LwWUvSUK8e1fi85EBBUdDZmenHknL/wMJ4BKIeKaNg19vpTHxArVzrM
zi4dITmp9dvsJQ5AjapoEVMRQR1CNKi0mmxePaeSIhxHi9r9grQmP5C7PwJ3
hsPcbwmSajc77BFVrqogoTILj4j8OPkUdJNmHBrYgXkgb2d77LXme6HgLI8Z
yQ9K3xqQ7qoTtn5vhQdsb0+9FI0QiVtXFWofn9OsLGZq710/Xrlwi0wzx+oQ
AktBNDiAXgHQP77lg7TonhrBU1hVwjdk69TywIyijo/QViFU3IA7imCKT1I0
nAxILQLFahS5R40WK9xOuvHNUlYPNG14wtj6nTo8UPvPjsLz/M3+dcOhxJ9/
c3uJtlvzEGrf3gDEYInH70wAQtlKr26nkRXXGqJaCSreTtG9ThEb34x/4BvU
lMhgumFCkAbeCFw7zBJzmOu+zcd0ZvC7xMzwy6I+PeDbRTLD87aVum5TKLam
TPGKWnkqZD1iaHXt9QKz1tV2iXpcHpa6cA4QXK+1Q7Zi3kgmzMvmRRAuD+Dr
N0R5gFOnbMTn3Uhws+lro6w5P6PtICUZv2pWwbRod6ebO3m/+E72VKaVW9Q8
Y2dZ/nWg7uLDM2Cx+QvVWBO9CGbNz/dAn3ekic6B/xF4P7D95iG+0WiOETBx
yMEpo6YcZDMk5qrMTsBhTXrFCzc7Im3rZhOUpxWMseIz6qNtICPjfoQlaUB8
FmljFSd8Ewl1AKORMuy3BTBytz21tf6olppnHsU+rXPpgOUo2tJGYPFbmbQp
oz/lwYgTEur95r2lJB0xmV6mbWdmWv1/GIf+15xAiDzysAedXcRHcYQugam6
D50gO+mhCfJ9lBFWhIMrp++CCdISe5ozOvXrCAEkC6nPEj+zf1NfjUa7krwN
l0CZDLNvizFpeyNJKBMCYPzQb/wLTvH+BmsI//eG2MVj6wXSEOn7+ozKiniD
K+GCuS8WSWgNbW9FLQYhbmJrJD1DRz7JuMY2gz+va0Vbypb65SLrn5+2SR+n
oDFtELshwcYfLalGa1gJKNei45KSHN4i8ucXvuwPjwteufxx/DRLtUdDAze5
LQjwpUtw0JhoOSMKixBTK1TEoBcAb3cPGhSaylQVxJLRE4Glij4zIyzK1Yrz
1FUKxChYvsZ5Iesrd7Omp3M9BUN8sPbygqPvOyrD8NiZMFBbd/VHtJfq74Lm
ME2NUlsKNT1wNAsDELvqQoWaVkiTV126mV92rxweoHJW9IXnoUDThLKkHxpm
TWJx8K+elXtiMxhYQmTmOQLT/Gz0goTaM3xDzJDEUvdAgC+Mqh2vRP8qvDF2
XFbHup0IyUzgy10eGl7W9HhEcK2XPs5Og4xNLwuXdfO2gui/X5bF+vsNyfpl
zc+mJvoKoH5Y5apwpLff/FsR+YxFoVSYKl0/UASUY6R0QVmRSpyGJ/Irv3d1
L+M1Bjn9AAw+AVq3yknoTM8kR3Lhv4Vy6pBbl0h+UO34nLNGrJ1elSa/K1Ve
sPkK4JGFUu4NCpaH69gEIggDN08WTf/LM30MCzGhIKUJFLK8txWfI86ix2op
rpUPTrIjeGWRyeM6ugNhwgUzfvZwJVDUS2UOwZ11EwBvJmikKlptDPEBrtTw
CGpfzzu3VvczCXH3cEwVIUAjos2sHmwwqtRRyGRS2aDxLO3BZ+mTk5cZQfDL
LG4o05l0lJ6TLG91+NUZw6STulya71YkAniMbYBpNf9XdDiWBH7YagU+rcBU
EaHitYJ0Ca9qVXNiqS+Idh8vgTIf2zsVo83qARoIyivnESuLhkDXQTkb4RUI
Iiph1r/cW28U4stGDd4fKF3KjI2SqMUhPbtc6YJyjfEf3vUSRdMDjMnHGAXg
vW7Rw6K8RJ923JDhZuXzMeFhT7sJQqtD/W/9EV6xzxU25I0Sm8GowNiPVsYn
2X7l73puCK5URAfzjOrABCdA8RebVRHK/X1eoeOhwO9fohcIf9+nkncqt7cx
esm4QdnbZnL7+QHJFzckLUPcd+sKyZPFsabGwytQ2QS2oIokEUDXgu4w5tHw
S4mCVA2KUszOkvRSlzjq5Ms+FdDPCWSey+fKwxn1A4IumjBUuYEmGzOe/A93
oi00/JjHACArSxpe406rzmpmFMy5rwzXC9XKjmuGoxa1XZM7f6jjFVWA/KJm
5+1P2cy7o1SE2Xm0jqG05bN3fN95ewlx+hH+jpdZtVzWHZZ/ZsZqdoTpakde
ae7mWO0J85FxpQIivMyAAWDLBruGPPpiyoPkSiW9zaBKQpuxiyH41ZotzkJ4
WwkkY6aX8HzNsFyZdGCYObcqgTQxswLKtohuM9mGNsb3yoFVGt/IjNJp8/r5
rzv/vrKbXFc/i6kiARqctLouFZbMXngysTo/uJ4SEYSvb+iwakVrhL8m68MH
tNw/oOXAeqcN/xBjeLaTHCBvqooE9SMk/bEN4kHrDwQ+2Yd+UECwu627wClt
IJbbaNQnSA6EDi06tVCsOPWtBf/ThsMEF17i7LBzoBhi+z7x66xrcVhHiQOD
H4ki40C5SCnDbMyhJxCLRy3kqu9s7o07ibhbGm0sAg7dGVH7mZyHKrHMr/+M
137U3HFXb8rxj3jYHzVrg9WWSTte7G7FASFQ1dS1kRQ8lGN4wTpM8fVBodhV
jrF8Z6wNHkf9+I5akTWKei/NSUu7IXtqI3vue7V61Ofip6iREcJnEsJk7mHw
+oNnlDi9Nkz0sRbkfObjGBXpZkSrPnqoZX4LzL68khyEMxGc8PGf7sA64BPa
RFYd2hJnPvc6zuosxZO6T0MBpq0jua8Fbl4lGlHQXt85NR6R19Pw44E+FRPO
v9wShaULcoyhYiJGcYK34Sdlduq1tsiQzrleCI7t5gTTthJ1ljzWpWQf4B2V
K/PcredrdqRQ4aPg5ENt4r4YtAkHbw8nET/Z1po+wk2JpQ1k06crKl4JmU0c
PkBU91ySGipkuSMK4+7CryPKxI4JBl0WWjxazWoHdCp06DefzCaME2wxF5Jr
X10pox9d1CYxQTT63FmQz9Vc95DLhlrwjavbCsHoH64tME2LV/Oha0bLKo5X
igfkxHkGDhSD18zjx/cOLAdcXBSlMEMVtjYqGAU+TME25Ss6MEGXFX4dxabo
AT7oLleiVoaW22Z8LwvpZ2UabgQBmQcWhKFLiOsc1XPXoPm9sWT8fBnFrLXg
NyJyRK+XK3aQQ+JiuCjI8fU4mFlwTK+43o2DqzkkYc75FEs1FkWLklIjyB8n
HzgcxzHn/dfgx7mpwjflk6NKUkmiGeFtM8M8xjZ27bDvITDUNkbNYvcbsVtq
e6MuTcfNkf0DNxM8UoTdb00dX2hyZeXu9bbM28f/5mrTF4fxGwnkWZW5rxg3
3+f/wvXQJXu/g0Sgh3QMuyvf8Si8U5OuBRS9w3zHM5hRkj200xf2quLGGfDA
Im0KSsCw2YQg92Fb0u4jHx5dWGeF/1UBsU2Jc1Vg8bVBJ1IY9Pho+xrKlziE
zpmD3XPMJuv+8Ebumnp8kIKQM2XLFukjXJqIQdyStp7RYdaTtYQgYfR9ezuS
ICp2BPCBJee1Y5VyG4TLhcR/0JrjAkxnPau3aA+FzZy9PKtktC4t83IxJJ98
rlY8kASXNyedaM82IX2mjJcpTy/aPuGtUs3qnpjqQrzSkZjR7wLpYTaV5kU6
4SZgUwyqTvzZICT8yGoWHIY6TzYf//6DdmRFJd+HZqbCfBW4lxiHqQiHOkE4
riRtDCeIHUDy7j3pjhPEOq8E4LcMCf824ibJUCBk5hC4MsTzvAoSz1LYOaWk
m8KcBO85c7uSIZaj/5l9tekVoYFKWuFgDskr5wmOempRg+W5CnxUvopOfkVt
fr4ByOP90Lolpa61YcTXH88Gv1AkWvGbO9+vviTGiEwDZs82Ey5HwHKTHym9
K599rQNfXGdm54tOxqHJ/096bMyJ++gWnZOAUlIRpaOKAuiBz0xSSIFlRjBy
8g0efNhhn1fhx40ZpoSmM3sv5JKGMyKiR/L0ZwEGP2q9Mp+NPXaXQ2tWN09h
NVHQoMYORPSm7OEfY3pTuxT4jKU7ul0XSmc+TqN85ZKUXS12hqf156la6kob
I//lE1cniURXDQ53NwSTqqZIcRI94ujOx2L44fSTxhxAjfgLg0gPeIetgq+R
aOYgWEUZzzCL23ZATHJonFswwDzPPJfEFBLNhTv7C2/Drtfhzw432tAp6xj/
VUB77IJlOwOFZEpC3HGnl4RfgZysk/XI132fvOqmriN5M/aSBeEhfi6Df0Wz
gPqGbLMLa5iZ12snCylKiziZeNpOjf48ia8ToEXFB28VNpfcujdY0NqNC3/n
OGvT2eVaHscWHYP3pULBPZt8vPRuXibtw6vnhTnK0mfoj4HT8QscrwbM4MMG
dlkN159TUcytA6sKeXjfy/EyYsyRB4i+taYXXDYl7CDx55Ouu+potSB24hKZ
hGPmAdjHb5Wsjog0RZBu0YCCQkLzR3BofAmUuXECAVr+K2S8qJPZVTElc9W9
VYkiQ8aPiSyoH9SI8FYfLgNxtChjRZH7LbII1LSlFkvjSMns+JQHT+GUOeIO
5vY6l4FvThNsKFzU4CBhS4q2En1o97xdGizd+tydoc5lVebRNzDByYy2kIlY
2/166dsykMvBnnMZQD/3PxZDZXfwbRLTwoQeIanpBGNYO8DUPV82r6XMIQ3H
8Kr5H9dUGCcroHD9xxtqJppZYIL6fuUM

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI1xsQufRtkPT8Jfs7n0skZHWyVOAB+GGiIoKc7kDycLYugEu8XET5XfCx6UsdC572+8GCk6TkQ15lV/3u7dQBuyVV2t+HDV9Y8R1KEYWf5mcuP+wLHsAq5d6rF0U2dU6d7/FD6hvglNhIngiHOTU945kQbOB+S52NFTAAMBojNy9KAQMbanYIsKoN1KQOoNr7c/IVDbePwI5uqIgrylBK+7bWqyQmZnINEVsaFJ7AuLF5Oc44xYBZbKuS0OHv2UKpCOMs65/9ZDRmxYIk/BOERLj0ygXLihgtWM20lVeVnXliltnlEDwJrLw0WxZuZkHlKEGrQOxPcP85LM1tDh0NF1dk7MFqa1n1eGA4h8lR2ogtD7Dcve3LfrOZ4D1Hwm4CGiIRsTcK5d7C0o7sWr0HwjS0J1ooCpEzAw99cwiHFcSXQb0tsR7q90u8mX1BPq/w1q3eXdDESVp4bqd9cEZY8+loFlJNr7J4sBUsE+aPbTo5wVUAvtkVeQxnaJNM7eMFq89pf8dRavAk2FGlCJ4VYkZG00Y0sMTthpViU3a4fDMIZ6NOMtAtRPWnP7du+ST6zvevmSLo9VSESMd8iQKrVjQpVcWqXdkd5ewmQ2cJukP9np62luSemdriPG0xy1/CMs77sCoUv7NNVD8XF3elqJUbDkWaa/FKjAbwJXD3oD9o203IEorZldbK9hkOiXBMMn/n5qYtJHL1d1uUG4nnXLF/3+4pBmU3OM4/jC/eDD/UKqVADHh7uJAU90tlespMwyDR6Q9GTIa3iC/7YbdLyu"
`endif
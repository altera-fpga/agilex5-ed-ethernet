//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QQGkUPzUaVjiJm5HO32o3VZGtuUZ3vTwxPRzHpvKfufy2lIQA1pqSLU3cyPW
QsqN1Tg/E3W2NP/n6tQfXbjxWQHRZsRQX2huQNpFjzRIxNM+1y3O/3k2qc6f
HTLAxfgpqqucWO8eXWwg9qpF/diT+E1Kmx79FJodw+nCZ6jYw8uGSlM1njk1
QlPNqS2vTW0nu5hiu2BL11akQXHg/np8GaV6W0xTdjRaBK+BiEPtMa1X2ao5
7/eMQwbL+HL2GARjfotCNSNE9XNmvmDq7b+6zX6EPcmRmEGJjwAOqlRUtV1c
LjBv3nnZ8fiRZMOZhm1XXEKHrBcTOa1JVChhwEfKjw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pd9yXAaQB2RKDSqKzxJmMCc5DZRIBsb+quS3ko5FjaVtwUBufMYRzmD09lKP
bkp5o+erdDu1NMaJJKsQVysoR2AyQIsax7VWImsLXdaYZd88BxKIWmVX0PS1
5yiAvcVgrPc2qtfX1KOPz6iK2uvFS/X+JUJh1gpQE9DDFqW+xuw2HkqZbu+t
anhIK2DX6GGHwuc0ttCSF87taRRfPe7Y4qbMPdTEdVSSCeR91Z4QgVWTsaed
VUzCOxfpxA5yud+D8foNghFR1guJlaea4FGe5V/u7YnbDJDECkYbSjvJcK3D
TPx7qIMI6tadfzd/Ujo1U1+49nisokFLMw9YYGaepg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n6GFiOsSevyPMt/2E77BC5TzcWCNHNmBG0iGZ9iz1rQZI9u4DDN6pItoqj7I
3/YN5mICeDcvry/K6sIFl0e0lyrL1Ujk+HIko1o8hIgxyvwRp7gwdwbLFaTH
rJ4dq3uuybVsCH/OBHU3QOJ3T6iEAcXhhDwvFdCS9pd7xk0zliYWQ+pmUiCQ
uR9NTGAvY+ix57HokA/B1uXypmnHtH1ABsofdvhuzkpQIOfeBnfA3reDwhKa
+p/W5gtKzJhelUVSTqnTuC4t1MQsFBbG0dBl8nJM6ZPpDHwCD4IptAzW7/C9
07ZELUU6oKefIvvxt4fkjhjvUnsI5a86hMVX2YXx7w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fxOmgvyD1qY4DRPnQVBGjkNrl6z/Cy2lELe2ypuaFKPHxxsUTuw58zYeO2is
C8JGAzT5wrNfzfmQly1I+k5grjV+dcb5dUvkLWbinGZgKbGywfpJhTPuCtfw
B4fDx7FBwFVmQ4yPGbWghIimEGH5w9ab1Mf8tVjQeQ+5PN+wP3AEyvadRDwi
WIDZGqe3bpMU7ugWEh07ShvQ0t4TCTidlxMtkHvpbqymdz4/ZXG5xlIKuQRs
ASdW24Oa7KkmVLdZFd+SpZlcg9Xx8alKUKQOczW2YHUDlOP/JERF7Finz/N9
hYsruwwQT074r5OgiiIQDUbUN0rHal/4c1NINQBDbg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P2T6WGaUERCHKPORKkPo4Kj2qUEJGPyqtznE6ijnRunVfueUMtlfCEswSviI
xjQwhk6gltGzUNC08JVG2UEtcblTAWlWmqXIO2miy569oP+POkPnwd+z2zuQ
p8HpKVc2lGyAWWmaQT/FxCFoAxQBUE70impu7Bqjm7A0EIRaUzM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Bqv1IbcrQvROa8pnlOP62iLyByY0wiCbICZsTbKi+0un0HX8VIJ8Uo/gaDUf
JE/0so45Uoj0OP4AMhxTTrdHjq/AnckDB3tsuRRQjAaAdrBrzaKSTSaLf/UG
UMVwDBoUCBesTBU040Guqw2+RUdLJD9tNkaeb1H3Tg096y4ZRFIUmhEqpz46
ENoe7dm/7sDp77P/1aiezdViPbsFFeXSqyCCO36GoxmUTiW/s/rK1znDiLK5
DPSRdON1A/xiBKaER2f8IAu35XeawTqsyZo+uAeXa5qwnloYe9BL8E/X2n5j
oNIwINjajZdAqQyBlgLj+9gDpHCiwbMTu+RCYra3HlKX1EsLpZ7f/bCU5plk
8Eo9hyPgcwhA+8GuE6XH6hjCjJDuHLG94m3evJqKp5hf+c0KDHKwLGJ4yXTR
ojnd9TBJaet5IeoZ9auwj5ujSqKY4FNcbAhwadVPq41DnlgugY6e34kQpCDR
LBtduFp6U0RiAijGd6t5xafWGY7IaWI6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m3XpNreuRZQzF3XwB3ifeHuf870/R+nX7wmPZXb9h8RCfGoe17CF4fuXEwic
Js9b3A3BDy9IIgmAjsGzwipQQdMwDnyZIGrnTSbdX7esCkt7kwrhOiJkhTuz
7TCDgdSz/ayr3cDyPSmSL2OXb7mNWXZMb9901R1/tuPQ8EB7U5E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B1PY1jv+jUhiTu9t+Wa+UfOwdr9Lq22ZHkwaoypKDz+KH/kU9YEyJEAUs2QI
DRcoqDRVEVC3FaU1npEE5IGhuvEkm4ne/F9KczI71+c+/7IAaCr39fJlUPDn
ozmeMBxVnfgM2z5E1yTpWBn5+loiDakslS7kx/2xFwMvlg6eg6w=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 90320)
`pragma protect data_block
10QciiFV1p1f9Ky3ZV834F2T/KOZirQc5/cwpOoIxg/5bjIg1hn7kbt2m/Ky
xFONusPTaRQuD/NjK8szg7HZGBW97Mi2yywTWr81/eYQcglzXXftUhna/Gox
bcP+6tJzBrtk4AcZ6j31PaywdpRXTg8fnia7hmdMCk5M0cbIFwqf6sEp0+I2
bd4jwkL9lMABNhHX9YNCnuXmqjgSWdT7Tk+b/fi5aegS+b+1eGElxDTKrJjl
cw8iJd+c7rpihKmz+WSrq4MpRB5aUcSGoShfI8+2W67YeFLRaupCdpww0mMc
poPxUsgnhUpG43oG7q/kLcaj65Bn6tiSi4EaWHA8QaeZeuXnF3PIhCCFOGFj
5xBT1tgaXtvFFRETGt1LE601IfGiEUAdu8WEHVebpg9QdwVF+XCJhuUMtbwC
XrezZg5TaCg16p9ORq0a7fvHfbKAmkrEHbAUdBp5R+NgmFhM6NWQwsdYtT3A
i82dL2AL1L9owxJoDbAplWJMh5py+G7zuNElCtRWaPdM5kP10lDjZ3WbRqQx
763xjhp+OfHjOvpsco82PweiXXUneJoxFzt+LEdm1u6wl0sK3htzZ+gzczK9
ZEJzfMc9Y4WB1uMzF3qqbn1T80FMSLjUZHKUwKQjQoLQvNIoXF7uTX4ZZ0ND
NzdNR2PmkLDwN+mo11tvD9jaiHTT5Hvm24QTEmSloHPVPISXiCPLUOUj16DN
PMjdI2U5LiarndNk/6GhrNDfF7nIZMeyt+3RwmDX0+pWDNUJfDDPL8lYwyhP
+obxtlGknqYtloJ7uVZjnLovA4gcR43zpYY62kDiYQ2SSp49GsVGJUIQM+Qe
IiGjrWDvM6XjgR+VL9Tn6+JvPcTlzF6vTMMKUFLP/9tXL6g+gwb0uaIcI6du
NwOb1HiZw6eMZY5ILpIx5PjGACldhzwdc0qbbKKATluiEkjCFCqKbY+1Fo2A
9Jp2KGo+XBHwgVLMKANYGxCHeUXjR/auqt5RxxtAkiFBjrrtpKNhWzjRJzf3
GmwWrmSHa+LjDCtgx7/QAEG7MiS79Abvu5QX2NB6Vc+TSCU1arOAvVlm8vs7
rm0EnLnUpUVtPIHE931Egs8oEz7F0ZRNxcgYScC/6R3i9eMfK+EdWJF1dnoi
EWQxgCZGtoHZTUxPwgy7XonYMnZX/atg6W+ZCJZFHSfyqtTYH2wArh+/PH1j
x7xQUJ509bPmrQdU3CoqhL3cVOsr5Ybfm7Y4GlCMBnHsQCGXvlfJX2QgbD21
J75ilc7aGcAQjuFAAzxPGRnzZnGFh5uzYV6B1BkPTjOD35Vv31DpObl6Na4P
DAM6R4kEckcFbvlzfdI201BiltSh6Q45orhXYBepS7zRjnJah4FuRuTAMI/w
1XAyhnS6JEq5p6A6CNB6fqa7TfAwxNo2tOjU8U7LypFxx7dhfTU4beMgIQpJ
ap1bl7TpI18PvaSlrHO5ehvvry4VIBkV4+zGlhZMCfHTeKJjrCgHf/tvYSHr
z64iJ9iyb5vSI2gj5PrUZYYaJtQncjmY4WzhB3Xw8Jl2tRXCFpKp9KPWjl3c
DNAWSNKh8P/D5DRKKfJ8t1LCz5I1pQcHBw7Z6CB5ZA0YalQoaUWEy+rwH3aH
yCPWtP6s7i03RwnlCj2C1oaXqIgUNO2d3v48jN+deY/ZzePhmdjFqC9oF6T+
KufkTDish6hvIH2lAUamTsIIuTpsMY6DgvE18e17+My1wslp5yoCGFnjdr85
tyD70XalyAoiAgPT2eXEyAKE3K5Jsj+RKfGiLxylH6TAqZv/L5Fkct11XNdH
mYEM7PUSWkDKjJor2JnVMNHTI3T8NByRQwM6tEFKmlE2A2xVd1JoZ51rPEW+
VN7LqVgncIZHZyTACdixJTfzp8Q/kkStDDPVFJErOasE+UGDAhy4JxqEpq5K
aHmqPT9W4xH6hqnyAvIQLtU9LC4yG6CIo0DVilJjc3DZtQSVOKV7QarCKW/W
6HeXB+DjRG0OFQ+lbsXIKRC2ENje/bXzNA5MFx46aiaaga5054pu3kxSjU4d
ScfCp9aYfgPBobDkZbsMHze0dStsQau5d1LWWjLNKlTVsSJ7GmCEt6sivAEd
xNBthD3JQYhTJopsHXgQ71AuHOAMDIxH56Z7yRqWvRmJDq8IU892OdV7KA0s
2N43BS3+d5LUB6y/Dtn7ICheYmEqN5Ek52f9GlEJ8GXHV+z8CI5+90pvTkE/
pw/0RlqSH2k8v1m19pulg8ucjBiU4Lvfz81qDN7ZJs+OpHJ3Q7emNLX9lHbb
emPW8Z/0lnitGr9WIicrpAbNw3Vo+YnfqQFXZQlHc2P5qZcPwlJM3IAzaSzh
GM4ru/j2RMlfifRvbEdH8YDHRQ0UANK6csYi7+9TowYu+QFnnmkJjDRMjJBO
snV3WndCwOzSUSgUCHscEvhN3+RvHpRuZgPwHx5GM1L7lY76epV845EG3mMb
KA1sRcEV3wbW5PoaSIz3IOdJWsGyoO/FwOEtkZkHPni38sZJi7gBbrQ/Jayw
dWp7foyPwBk6aTn9M2CH/kCUW26YUeUHUulvOoe0Bt2WN6+Mnup6XIwsUXnS
kgTkEosrBmYUPq9hd2zi1iCxD5J2E0Fb8qy67GDCKy5LzhFX2JUxmLZRfJoy
lRxLOrjRK4ryZs7gXrtf8/wr/jyKzr3gQk85dkAmNcRzTWmBMPk3MtyHthQy
G3/5iMny3A7kcIm/zh5+05qRFiGTCSLzFmvGuLlBaMnF6aJgw8jFjMkyoidt
PnZQAyWYhP4BN7H/5Y0ZaFvjkmt3ULQe65aZCWJ3PNTAUy54QSNxyCgvKiK3
V7dHDpd1lt8IrfozBuO/V4XbmQ5dnYXfHRLbzFqZZAFnb8TuGjfqmXld8uxe
n+89jLW1QoC4Xt3gzWrtcV0WBOS7/8LfjvwhTohIXOzZYSruTNoQbGxwPmoI
5eTlsiKokhemxd7P6JJIwn/a4gwBYwEzQKip3G6pn4SADiyrzjXS/hRUGLeN
dwyDGSLg247oZ2AVohzop67c4edrSiZhY6V6BKjlHo+nQCaYla2Ns4McZOy4
DPCr/EPR4C9OZddFi4qQ5eGvx3M6VrIDGqMy4UaJMTj+kcssIvoblJOUIbtX
UzSu7Wq3pyTsG7Uw+Y+z83vn1VcG/KowXCO2T65l4l86+jp0yiUqGYL3w1tr
YXcgRNvEWk0LFBXQPj1l/MJLIO4GIG03ev7JhfNXRHFgf5uHxL8np0NwFFcp
tYh3u5AGetYz36BM9913mDN7P9kQHgemk05EYzd/Pn2K17xfoAGXUQg4oqZj
l4m6fUsUEaP79IYEna9yfWwd1oGRInpUxrN1sXvW1wD8NzecIL8oD4eoKGsT
K+9bXspO8jMe5fBhgc9PShuJ4zvAn+kZ2Ow1VhlujJJlSm7qBLetGNRm0UAy
zaA8gafhlh1gF3bpQwDk5RWcVg6A9MSKcbjDi6DT5ngpzhMEmxzI8EZP6d06
zlOWaRhMk3R/gW8Zs7vfaBvyIOhD2dnYreWI57D0lZoC97DSEFWfx6L2mm+t
P29AGQ+og0CxXy6c2+FHwqV5JyN8QhFxexcxZ8FKvoFb5e0bIasAcUHMyCtT
tXoMDq47ArprHuk4733sYxumTlBZiek/aJUhPTVEDJ8Dr1W/ok/coSJoVtAw
Sr2jDiqXnPmsdMf/JYTOyl1/EibOh5GdlHbFNEMAcwhllapzDD2k3aC1kuVC
3H/JuGpYD+10rkWwNM5n1cdvsuhKKL43fXz3jI3rmcXiAZVbGMlGyPjeEcyw
ZgA32qJPaGURljbcGcoWd9qlB0e/J32gQhTTFLbku0vaK0Nx+ae4KY45XaFr
Cw0nDK0bU0BEHMSjpaxOeeyamv2ghihjvonleKLcCO6ixQBzS+2wpAHy+o35
NMPhl2dZJDtySJnMWVR/2lgrXR/FH64O3AlpJ0+mjb2MpW24wjZrGwojfC+t
D5CeaqBgQDuFYA5VYoMaXdMliwl+4dnC6h6aXfLYv1Ru0LWXCpkmyFR6U4dh
6qD/wkKlnEW9JHNXlBwGV7y/KvQdX0a7PlCAgEV6BE0xNfDmdf6tm4+vsGyH
5khRr4JWzJp5FkuTzNrU9ExpoyH580KMLfzFqw7fq7zqrTnofhQCgZ9k16YF
Cw44bLFOhgH9nVRmncz4hKDcRHa/vbFFUtVTTDj+WuXPF06hyg+IUtWhIznw
0pYLvA65ozub9XZMo2l0reEhBlVbfVZUSYIS678+x70lKDvRtST+1nPnYx+5
sc/+ES04ObJ6PxXHtuqtNqEsaKCLMYYqHqW+fGFi2K5cqfSjDJYOxAr/A7cV
4WTEopRAHPbO3ah6oH+zScg3YZUvn5eLDPeLeEi4RYqUWvFWiBASu9BXk0E+
c/23P1/2JCmlML1y6zjeP8jO7bN9ZeXe1b8ptmraUgWK9e/60x/oKvvqJIy9
8E3ecv0IjKkukl/VrlRpDIsTqXHrvtSDPMKVAa0OM5ZMf7SQs68v5lxaI7Pn
+/v6a0U7Begv14e45fWYgAP6r1QOx2+hKhUYfElbeHYGAjTx6YaJKuQGO7X0
uHF7hXzIvzD50IK/v1/YpddLJJTsQKJ02/93XQS0RXurgNDYi5rq9wy8GzAd
MUXBsxxTFpIx1ruLzTPrJMMtXW3Q0s4LGVZAcvEJayMp42f2CaCg0aadEe6h
YJEwTYijqKF2QPJxprZ37Ch1u2/zGbeLWoxZ+bGNXan7I6RpLrY9MYAy5RO6
z5SIcCSPmUU9SyjLW+4LhElHXm16+YlEEO/+t6mcaCMoN/GHfquEEhKBra/W
vQOu+uSE54qeoE2u+baiOQ4PcewMcJ7go9v9ndYScQxMHsQgYUjhA+tDw7hx
yJ3sTF9eouK5XGZ/ALOUPM/k4+jDVPiITGtRS3AqnopITRZxh/eOvTWtjR7W
wqrzAYvgH5i56rwbb+FjmxGutzIn8KgSHqhvh7Ig8/fscKYU1k9/VIkToDCo
jRrAwema+Hi3pCwU0Nwepm8GIJPOdcGtCuKb0HDCNG+ln+xaHAjNg75DIdEG
dTG+c73PLRMqE4prcU4Gw5EKv4PSNzodrLPE50op82G9M6jZmMgrBVCICz0X
7hxgeAGBtWb6xs/3ME2fgLjipilPvQac6pZxIx1j5FGEmCbZiLqKXBpUEpUo
Au9b640AvUhdYvhtGUNwevHYhsvmfMgRjitYmrk0RvjoysgP81IX/o4mRLUU
3IA/EXnCHivChTxZY+y7EipZb3xpR9uOTteybYQm4FG4dMXiRPWsil+cmmQ1
jJVO80ia92dNpro42wqkCI4IKmqufET4v14dCT/91MVe9zeiLZ65wIjJ0uhf
ZC9/ZSS66WEaTG4EklO/VnPoPaZjDP22TcTIJuGhGpkCXWlrhTn2exi/eC9K
esrQlbIOqAdZTn0K64Qz+5o4IZ4XZOobTFQbv4UmGh1KxPYQ/mk5njFrzOP/
M4PxjpXM/6kBpfFudn8iuxqVMh354B2wQBOePNVyvVlgn1iQDM1CYXpPlT1o
OSPbDHMtvhLXAq5j1NU7f11J2h+lyZvKTTeKt7h3cT3exvT3ZSIImQ+6aHHz
ZEsYDczeIgOq3CT8e5WGiZrZEV/qtP+FXyjYngF6us8rf8kNzHw4thY2O6LL
A8AAB7DPmBI4LjUN8CfItK1fy1JGmy7CSZyV3KjRvo6Qwrh2vRSycANGCuko
G/8VI6WxHijJWL82lnHk7j5UuRXbIqqz3LAWyUx4YL4ng1EIVAjjaO/1YP8/
7PL3M7aY4WlgQlXcL8kNWPlb6YPUvgQ1V6G+3s5ttaBnhMtEcd96HnqAwkXs
TZkI3crmqkP5tWCcyzxv7YAlC2vAe0qQzuylnEaWhTMnsuuW6zrtrU/lxZaj
jc+5sEzImDcof8TwEmfo6dUpR8bUWDimHD1EgVlUiBdBYuSph7S10e9Lg6jd
2aZv5xUG2PMiy8XO/aCqfTXNOcCE+RyhmkPuEh3U0TNCJI87qtgeoIqdae0N
kqVIoFGnsDKbQRbPqVgTn4BeyRyT0Hodoo59miRg281/GMnoDNrWFZQeKHbv
o6F9Krtxn5t1D05HOwC7jI77YKAZ6RMWv/HCxd/TGTn+dNv/bHOGqF0nbJuJ
ccEx5nOeSC1w5Et9tb4KLXagwxuI+HClQtAnxKcgwKSq1C2Xg7xyc2KlL0Oj
aVhARtMhYWdy9S8eWclT9aGolGyTACWBqDIX/UMpsKsshB4nxKi/pIIzmAHN
aKluqVE3fkVY+JB/zpZ6wmcSUCo7ZM6a4UhNPX3sif09K8/vRcclpz7PQNAu
k0KsuVWfbQsqrjFeuic3CF1788xoJgQ9NEVLW2vZ518YdAvSbtO5E6D1cNdW
RQ8DRGzPtaGtHvsKzTHWruRKsMesMl5qOs+zeF2XXO9F7DGpWjTv9E86Zw9F
Qa3ZNPVk8moj4Ok151QZoSvnJRR7peNHY2DWBPV1N272BC3PHIAGLVU3r1jc
qPnjk4+JZ9mhMsvspJwJFNRT2svB/sgcnxvUs+7W+B3W50OfzmzHyRUVheoj
MtY5YTyKXYjQQ1ZsvMQe6RgZFjkdCt3AuWJ0aA61QV9fzgTBRcrMNkyLSd/8
Hg8BDUIee6zVZsYmqs0ek27tiPxnMesLtgwHXx/0aY29yw4rRXarDRTuvDP0
FvqbUsnTCF/jNW8WTKQ/ewIOC6eADbmnoO2rG4UxqT4CzzoC2vb8zL/ta8FW
XnN2UpStzs2eFO7q5rX2gd+PLG7SVHdVyooSTVaz/eCMx73qHTLenTMQAmkk
SKWjLwLFAoGmxdr3B4S82sA5HIXpk8Vh+V+pnJnEzMK5FG47iFtq1Ot/VJHL
L0Hk8GdEGjHIGbHNiZ/x8mylqU/kv2vOii8CjeSCW9iZ4v0y6sUxYiL/GHo4
gZZctkKni+44dU5CHyMwYqrJAW0TlTZAR6fbj3TSmAygFFUn7jHNAtqv0zcu
/f+X+UrCDPw4sRN4wwrHwXMqE0HdFdbFdHVs3VJxf9ztmgcui0T4etKoOlHy
54OJnBHKlDwuPk+shfy5obe6r2JQdKQ0yRWh0iyYg+VHulGQitb/97mDe69/
/dczl7abo92Z4peIRsyBYLqdtqEqG2e7knmyzD3MO1nvTCL7/qqd1snjs/C0
V5+H7+1XuUb0UML2CUpTLNyRCz+vgqp1bcTMTtS/AYOqy6AKJVxfpGH3rcPP
xZEaO2DdLqAL6THr8wmvYyfuUs0LyNpZqWLeDcuGjNqJaOgEF5kMgJnYrm7M
o0gn9M/GWQL3tRP+MNDgzESKNUOFEzfeCtDLhd+ws2Sa1nbMWM6qGdRaJWmY
PTO6FfIWv1U4DGpOdc7kaWuEfzkVZX+tpQd+IkAkCHFe9zyvySBH6VAiaroT
AEANftyvoXzfRKGeaKCqCY0CGoKkYYvmXJjjc8m6jMQ0JzGscP+mbxgE9yG2
pp2G8lpm8uKNtoaEl19RLbok+tqAD00xUzbpIQyqJEY/lywlQFGVzW5+G4yf
cYthFPOUcbNHlhVgo4gitm8b9VbXLSp2ug2n7TN5XH66CYLFamft+i/wtEuW
i6/8Wp/4jxigHCELTyh3OaU/vSVqdI0zQNz5pePmX+fMs69E0U+dLZZV+76p
SFxlTWGd/jK+Po2G7+ljNbXNQO8ifjG3iNNiT0v08MED3mQrMzTunaHuaqIT
PBcAsv17XKd1oG9AABqBHt2wqbWwuVt4wW40icl7lOsyu3CmnRxoFl1souRD
FfpMmIoqkZyfVQPn/m2TA6SL/DcmOrQatvlDNlt1DpeNcCrTehsGFLt1n3Pk
x9lPGF73Pbmjg2pFgbIVAvfGduqWYZBxVWOG9tdJJ/VWeYFEucnIiZfJf3xW
EbBK5/OtGqMNr41btwVCACfR+qXz7DiZ0D94QW87d3e3nUzoKcSEbv94BZsu
jJ5aii6TyVHL73tZDr0baNnfOvgnpDmZwYPAHFanfCYPsio/rY0Okz4FdSRU
NYuJ1HR0JatUbn5kXaNsoEEBYdKcLvPR/UAE+TrYNaHk1kTeT92C6/RpFEtw
yxd8a5sF3uF7gkBibnWNJELymbXVbp21sYCSM6RIBWgWvH5H5/dWpANcn450
fy4LlVaW0uoQXWACyiD5M/cWspJmf56LnUI0buxMRQmehPR7N3KR8k4ldKtV
frRDqt8j2HJ32dpa2klKj91DriTxgJ0riJctB+knFxDTbc+tYKXIIIW4FRXu
CxNOm2CrkL+xOuF2JcZ03xO2hZavfXIiLGPMdsWZKYhBY3G2rlf/IraL9PiD
xzhxz3FgZVz++nB3gPzd2waIkp71v/mwTF0eTKpbSal+J1aNiintzN8SRCCB
tRlS3s9iJZhOFop0s3VLHwGrViGbYnCG5Ry+9pN57H9ojhcpJek+UdulHLL9
AKdeUW6XI2VPMwqCr3L1nqMCuoeAM/REeO//wzYLiVnBjeAlKgRFFJX+j7Ry
wG0+il9HQWP0CprIXP30+LH7vRdbudFrYjZgrcwRub8GnnmLdX0Y/+HiJjXO
9IGDkaRZXP5eNCFi0P7w5GHRxkMFSz/5+INL6zQVTPmLoQDXpG9eIl7Pn7ZK
VIYNxRKGWQXXPlKq1yyOaphNvTA5MXuHo6+vFgUGVL//F8/gHGPBSzqu4UAt
/pq1CYGG7Fz+eB9vNxTXwfFtz52Kx3KQBwt0uPSzL0J8rVSDc3mViIlyYQS1
149UaE2Q1g+tzXfzWOilWi+2ijqVB2RNiDgV0gKfvB847eIZNsnCdrgN/O/H
eb1mjQ9FpggDYVQ6KUSGCCloQd2+1zr0f+cD2ohOHoIMJ0EsQnVH9T5zx4PY
V40HmvfxVBwFeHre5OVC5djJmQ6Be3qABF8AAhPRU4WZzdzrafD6y7XjypSw
uBi3Vka464iIuzbYCh5wz5UC2bkZ+cRMItitexuL3QR7Rqacl++77qpXI9i1
ayAQJAwFPfbHXlEWoUQuD+ZVrtzKjnexqVwGNREbtXBrfFstyf0aBEaRD9Qc
0KEiIFZaDXe73553tAT+K0GG41IrzcQAoMKXrdazkZ+Hlc42SW01l2mVXpI5
EnpC1qfvhzw70XqY95GO5uKmwwPIgkeGoCg0HtFDhVLFnwe3ZxU/c2Yug0Zk
j/WKcmfsRNiFi3OTGqryGhovchckwKxamkvfkyh7j92MlAoxmN0AZjFw7YWL
aC7JBFoLe87Bm9FAeyhHoPhHGXXuzBRRUs08PmD0sNyNUoKYZ5QknEIgShO6
0/79J42smswHo12/wrxZ7jLne/MtHar9aVBidWXG8uouhtGJU4CuCpSAakvP
/ywuXWFlqdwK+/k18Xc5mBQ7DUrLYeSgtw8/A6HS7raUzySF+mMoIJWYRkc7
yfvA3qgbIowakiTCpVMtSS8EUie8gjp9CSmOcXclFEys8UKUnCaeI6Uff7C9
/bYX4DRv27TSZcuImJOPfY32V6xtMRNmhy03/oZYBcV1YGrHcZ33Vclbt0kU
fM5c3n9YZeLUQ18gSgIMN/dte1rBA5YdEA6aLxz2SLh2hRDGzwwm+Sj2Hbin
Q3leiRrdXQf0qUwQtcK2bGHjONbeVsoqe9xHN+iDOgl5V5p6aY8+zICXOhLu
qPlizor2aTFOEbXoIS9erDN+NJ+ZyGWD5yOkQCCP7H569CLr1OG66NyXCHXI
V3HJWMP30Xw4psR/D7vmtOJ2gYeHsRHjmxDBP++IDgZur6XBCTX/dbVjrTXL
5/O3xAVciKFdgcb8lvH9LqhjgOBuKGmrmfunlnUoaNZgf2y/pTgsPMKVVUOV
hBm7Ws7s5x/OxuGqF+eijBkWCPzNKk6NwGeMJiy1lJp3OCn6l3KANXPdVp5L
GSXRqPF7LUDrSdcGnylQzoYCypVIbMIiq+WIZwq7kPRKqqBUQhMMvQqqPnaz
9P7g0JSUCIsU0ICHeMubRcifkMdv6M2gA5+SYjtwP+Bhpt+GtARf+cQx2Joq
vMtm4Iea4yRPOgsT6VPg32m/Z/KwRN7u5jKDYkaLo1lAHW+dB9eFrnOpq1Sh
/r4IGP+t4tLlxNdD+GGHFvrUe66No4w5ZwQWny8z/pEOVZYXXh+IdVLrzUh2
bHOyaFVAcXDF2CrbLzFC6k1Sfcv6MD8se2AH3x4t8xZS/pGxCpG1aWIs2sGO
5CGHQrzr7IQcSvhXOPVbS1wxKC2l+tRhUjTn0Wbht4LfgQprSqNEX6hBqnds
4UUkRQNHRmdOKBb+Il7Ku9NjqJWDwbIz9GPIEePmy6/sMOSohqKJpvdNWhXW
fispll0Q9d0z8t6WodVCHBIq7ujIYxIcXvIqUOobzVv7MJUl+CR1g3UXzBkP
gx/h2aFzlMnhtsiWE/+14hm5v+VTaYyU/rMWf3xCeYHltI4BDHQ9/qN1G/Bb
8gw0wa9Mbjd4mol1NDcTA+hV5wzeM9RaY3ji6CB00wyOYJ+e2qQdbl2nltpV
f9+PSMtOc/r35TqYEqNPi1RKXzQPw5SgMt0qmbqwfnhvWxOYIuyfGE2W8uTq
KIA+PhJaL7M7+UktOfWe1p1bvc8sKbdZCAOQeldhSCJQCTwps3TWgs5o2NQM
7BUe15i86vb4RkWuznJqFyEAcPEvC2ca2teNbmQHwqsUvlS7Ys5g2tARLRiz
PAerSnj+W3Ud6mUmTOgVoZS0AzTYh433y1D3P9YaW5h2uSsco4orHmQv2AwW
nKz5MBPfamOtW+WZ8U7q3rjajqKwQZ6mK87KwOwV/QGkrbKKDEKGrpytx2Gl
5Hx/X2ZpzcWFoS4+Wr1TdDdH/v3akKx101WxBZn59c3Xazy4Y0+HV7sUz8qJ
7/davebfQWyvYH/NZWLpHXJGgr2C8OipwKvOOt0Yt1NOygwnHJzH/iozO22R
r7204t88MTl8pgEl5h+0IDju2UGkTEvGpWxgFDz59XKW48KfGQwVWC++17bh
mzbvxF4611eZuL+KGwEbBlCIJXflelwO+ef1tjVhbRlmErKhK2V8gnp1/qpp
w7/65ZWABIRqy5Y3LvC6m0IxG/8lO73ZL9z5XTWuBJjAUOcIHAk3UiwxcfXI
6hJbOXzqVUhMYb5tMSgDpaLyD2mVDK7ka2F2O68v/k0bFx10WQM8IuH7KvPu
cc8f/EFQmbpZFJ9TvmJMlCNnh4PeskVuauIKn6Gq12eJp2dg40xfTEnzv1oV
N1g80yynlS83HpYTXgjJluWHFHW+MBto7Fu95FJode5M4fc6UP+MkKlCTWYe
tYM98kdzTMqtyf+AM3s/rifT/0pbBaozsNWWGfAPuEV+Ip+147N796dgFgPS
T8P18ZfDygTgTSbwoctlyblcRnDKICouaBeFlW5R0yL2dW7V0BGrACNRaQdG
XS0TIsajljdlKDTEHTG5BbAYICyA3/o2oxe6DoqNdPsAffmIqg3FVYTTiBMv
f37B3fAVK0pah9gWGCgUY8L9pwnsOoxp8bxC6et0lb1uTiykR2fA3RUtp+K2
tCyAuXaHW4KBVmNuPi5QGDm1P/mfy3xiaY5Vav/pdnIu2RbyMB5uHeTuqraV
2he6XNgK6mu4qTd4Y+wBTMh+NrcvikOvbweLytWEdJ/N1W26GS7kCpOMqcR9
VkEohYSQMZ7xx+VigRVoGG93ULUSjyROTzRIhLqq3qtHWVuADQtoRK8u2pfY
qLhls+pKtPl6ZXSI7VgljZ+Nb4+jDb5egwj62/OBZAJLEtMFkrbLvVwHEQjl
frSYtLXHxuDK536lBg+aFXvuwpMjF1keYuCPRQzYqlqzFOj5QvUJ0NVdNA1S
QMvSDD3Ndk31oF3kgcERpDW7KxOD+L/DPzTnGdQvfCxQw3uJYCDINvSPjOsa
o1Y4ag65kEKnLJdVGnzZOSCFYjcI6eFbL5sb5ParxlobH/5oP1EHO/z/oCNV
SOJax53PjOAN+0HrC1KcD4GlrMskk3KXfvxqLu1pICsuXic09YMeKp0786EW
5H3EQGbHZzRo753OUjj3WwsJYyHjRVSrHUKJvANPvuwbz1cdzcFpdaH3MD7o
pBXahkEAlxW8qx2AGZIQu4cpEGSItz8GBaqNRaP/4T4RvV6ZwD1A07oACUyB
cbYEzNo5isuIpeCPM5Umdt0U8vHWBY7uOl6bGyDXGPmj2ZpjFgn6Rei9gS+u
zc5Q9qpIfy9Tfdkhq9SWnK4XLVlPcThHw/odsgPhBh3U+J/rkQfp1jn+BHK7
tonbExRYyAA1xQF8Dt9Pcj/0jlEHbc4rC1GY7nyEjV7VFpKDc54b1iTtaxFT
YerwCdVVPy7jWZAhbwMDbZZaovDFuFiJevVfi3bfh2/sSr4OvmVBgAW1ZhMO
wM1oGwcG8rAofEhCpH7HPI16KlfB0ipTmpwQBnLa2+o9mSoH5VQj3P/zj3Um
FUeXmgf4yjipC9mLen9Hh9Jmh2MpjygSetU9NOrmGXCtkghOOOdC+of8Qatq
bnbxTaspXJMY77L3ixV2pWhxjHSyYEiPdxU7C/+OlYWlYugcJ6HLFISCOVsy
yOBl762iLIKp4QsRSXxQrB6LauuA/RnN2Q3RHAZbbdjQiWAYHnjXN6LUqTAy
HRZ4x+CYQ3nvK9QqHFC1sN88wMB9AlSVfjwzY0wQSnbCFHx/N4xrXSx4uW7C
FjI1KfV+2cqLaukXTekkrwexFug5FSR3TO2cDRJIbQYox+tXzKbsKHLGczaN
/CHpvo7yAipXxt9qUXrsD1lCdXhRJs3viQk0xcUeE2/bwFNPH3ek1VH6296e
XU48LRjHA4Cyp2y+k+P9jTe8jesNN32PzHjVCG8LHPbrARFvy4go3AM9dhMz
SDZM8ibeaWtlsFFX42x1QFoOJ/TPlQOIbEuanp+9cjJns0lbZCFOB1ge/HWI
u/FOTILlgv5nvg+6S99Oo3t92jISl353doFc+RteVQtNOQ2bwmiUsEikUi3M
1YpIVkCFugSNgTOHFF5jsRv6KNekxAXL7SNvlUztEg0r+vysN3gUtchn/Vdo
i5vTHRGEt2iBQApDjHnwnTU+SNjkqhUnUFG2Uv7ITSXMKUoPyMVn+bL4fIWC
2b24MUXlx8E8kQ6v5woKU7a7sAErqEif/ds5v8cwjnOsxo2BXQC+BlVR9lxk
a5OXVjCGGj7c2TaAbhtDQ32lEKDziGW9IXdfmAFrHqoFOg+Uxn9b5AGhXD3w
cLkV1nRpteiSSPZkVgc7NzYvLLgPisHRrihbMA2dc7Hy95S/dXWNuN3HcWcB
MNs75Smw1DJEHNAY61LvAXjxEunJ0XmeLVYyBnNSwEIplxEsJEafJtZo95Ul
nlltmxP4rref+Gqf/H+D3s5QfrLpooIyEzoLw34fDrgczKHcJBMzonJIOfio
xnePcoMSk0cN6TCkUt92EHwSFE69xfqssnKQOBbTgBD1678Go/q/8SqtV0Zp
bXzSTlDWdh0sqQMw6wGl9xfHEf5PlE1utGpW1WkV+k6aejKBHqYvGzWxgxJI
LKxOjG958w6/LS3C9pqhylVQ+/uL4XQSFpXBWn5MzqJs8vdqrYHUmdvaEORg
vtby1xzMxS1da0pO3Xnhc3YjP+eIN5q1w2y1qToeSEH4AagsMXabT9gcymLo
5Jr+mXtfaqZqRZ7dcLVjf7yIg+FPWnjQ1XK0PBqDJYBsMNy+j+o4u6s/O/5a
wu8o15rHRMYU9WzZ+A3j1fVkvXsDfVzJYJxtDeBTgHlXAB1+eLzzoo9hpjEy
p3a0WK0bQPt6U6vJHMdGeSgBPEvw1uovOP5YYav2Vh2rRuzlrvYQVzALmEsq
Ze6Wav19JENO/y8K9T1q5UFOQojsFfrC7J08413MqhkIoMIrDgOMsQIi6gGv
w6rrV+tfLh668xZb19bOIZRRF6Nae9CoL64bkHD4d/PJod4C/ednKoAWiKj4
DVtzZkrdnrGxgBoFeVqWFdjSZDPaEozSsXkSRRnuI44Qr//ls7uXRPPIM0dt
02YaJDNP4Nk+i8Fh8kXlKgWxRNgxCGtJlUTF1cpbdBRJHJ8awVgvs2JTCFUY
AP47zP37pWlME0l0EyQKBEP89Cek9VNx3lrhND7CZXGHKqT+P+AJMJ1R2Akl
3raWEfjmQ5jyt+l38+o+1Q68yaecJNtIckeDu9Bm+QH10vdLsCi1wBmvshTE
fY2nB2GXnbMCV9j0BDdWZw/epnZWeNwLwEsW+eTUFQnVPtoDyHmTRlre1E+Q
ebxQcPCV1ew0Cgbm8eZq1L70p8JWtzjkGCcaQ3vLVr5sND2d59V1gHrhfzgt
lV3pwHMB8MD9cdTWTZ7jTb1PUaqnP8AAt/xi1zd3zLa6PIcFQ8sThlSkjFwT
CafcXBKpnJJMCeyLpJ+yhIHHfdRXfHlrJMz3fMB16h5u7AeGjOCBOom+2NPX
BwJkuN8L5LuiMs0nVUI6dShS7pulwNxLxl1+KJe3EC9mLaZfzFCEDdkhvgTW
NnaLT7pbrjIfJ2pZDijPgPNl+7aXKoG5Qrxa0/ryvTumY8hd9l3qdsb94tng
igoZqX9zZ31qfjBtk3AqLql7eb7Skpf+gFtc4pVTH5Gk4eSbCsd/j/meUUv4
ngL3O7sG5FGpDb+qZJOmM47gjy42G8ftStRRLBfRbtRqLqIJwabem+D0FkTa
iLlVulVOogD2bY4qPlZB5Og9N+3tnMlBqB1APmtOnIwVmKq9c9UwhAf0adSp
F17ILK6bZv3nOpF2zfjX5ZU/NAHPi8FiV6HuEuoU/COZoIt1qD7uFYlhYkgT
FYZzNGJROnsbC9+au/8eVx7g0g6CE5MBXAtul8dSEoZKdg6KsLjUEhfwdhrR
M03rSn2WsCjCFrQKVrstUK7Jzzj9Lz3ZflfENn+hJdF17U4u7M52hQRI9pEn
njzM9TwtXuMt2s+z9YHXvut78MwulvoORenMg9VuCJgklKF1h6lCsuP2UYU6
7SiYoWVHU2W02ufdeWL1Q2R/ZoEtLI3ejEwnyqABPwRusRTzEdPjW3dgyvhc
YIKocBcxFkvoomnkKDCAg8ruCxs4RlAUpvwEpnree6IhI1FiHggmU8Jcy7R3
LN0q3frPBD3N8be+Wyb8Ar50ipMd0J4o+LQrmLM1JqwCy5xODFNnX4lpTkPj
LihcwYbVEwfik0VUL9ZQkRQhWmrn8bMN7wRtY6T0Yhnchex68qRf3oFzjViy
VPm0O2aWT1scmAVNFFC5bZ3DXa3P2+3zxkdERQ59luMoUtu+Q2eUetuSdSBU
7QASthXZiegHgv8Gf934ok2Mzt5xVWUwzUV9md4j+40v4Zz4/gsdY+zsY+Oz
Sc84ccY4OlahRd7PxG1NL9XHa2UVzTxy8xlOLxSL9EI3nfosy2DoQddtpayl
pJSRFRrcO47NpBt5tOocasLsOjuW/TZaHRU1tLSoaMfCOWK0WpwxM9/h6PXp
XJroznwV9s5jwwpg4zBalv+Gw6X9IRvNmAF55ovGI4dIjLwTTG2UNjrNGmf+
NbSDKk9MHlZmWPfm7ALUeiYDmwmsgCeyTpKTdJ3zXGUZBoC8ONwzW2RUReCW
v3rrlJVv32A7OB8VXEnPwYYxpHXoB0icsR3VFC8KgT6VbBtBszCBqGNps2UF
Yb81DI3NlDfplKB86U0u4HEJWQWvixjI/x2W43NV2Kxq3DBz23SCNuebpyAx
xj0ErDG3TfptpZCYFkZSSNEZPdq6spIUVoCtzWhKGyjfOjIOA1EveU/wbGiz
5tKvcmz9j/d68fujcE3z7rki2IgCx93b3DSrLDPqJDHfRXnVkDR0twxejYGh
NhSbKQjIj6U2WwDQsWXZpxDBPa8gR44JveV/mcRjTmSwRnYHQtyHBkH/P1eh
uexub/B5EbqWl+oRmwewbUtdZPswvW2ePJmaHtPIAMfY3xaj0bSEElI1dvWT
4kXgTThF9pBXhte8cIOo02ABitG/PJioixkEJbIZGYhUeuZZsY+A/KPKSB9+
X1nc7PmsVR5io+CG248D2bZE5TnmAgmJ8i8n2EWyAa4KKvAsOHYnHQrMYVoo
cXwjG+ctbAPk8df3I3PbJT2zcqAJjwhm6WnHFKaeXd+vGQSOVf5ikm8miMBk
gHx6w9U7hokWyVcpG87per6e7QKIzlwvOSJ00NT8tVboarWsQ4jFE5GWwJHe
5eaXYVcp2EZ3UUezaY7SzXpjR1niTZ1R/bo/Lbi0x3YQXY7WMtheW7r45zo2
5HEj3CWpUFplgZxVhLP5iqpYomnBSLbvu6Aq/fTON2BBWjy+8W0yDbJ/Pf+w
MUJRSYKRlb1ZOn/r1WprbKqETuQYyOzET/6huV9UogoYG8ZmTsdAU5LDp16j
Eyx2yud8IWjeGEFGU3JYNan9MFzC9tmjOSDiDrcRYzdJP2KZEMRni09o3QUv
qjvx/QJ1GJ45EV4mwe1P7hRJROtI42Dg/L78n9iXqBxCdlV1OqvFgVOS2PA4
6Tc0N+tHGnY2QmZR84L37cBrcEvFQCthQrlWGI9ZlZYlFjI7KTYRIWUj6UPy
ySx0muLlRSYk7klW8cyplfjoh9851oME4Q4WfOP07sfcBjye0BD/W1TjwSmh
slqXlyJ6lOmjNYQNFarI0xms/XVzQOrGQOzFEvH4h/a3WYnoC60GRL4tobx8
tpWO6qozzBvUOxpfyixMnBwBj+NNEzqYlsWjqKqkuMg0xS7V9lCP8RmvOuyR
e/ccMGHj98a+QhNCOiMUM6FXHeBiBHn4AquFb9Rv/0BZvwtsuqQDDOJj0TH/
87s2wUNcDvU8aVbncvxieuFS2LcZJ9+ig1+N3fKRtIJmHhc9Qy/TNlmtvxUd
PMg/KmoqwyAsvlofEo/w1PepzE/YW+RTBUQ7F1PQ5PjGnK2C1o5a02sf/iwi
Ie9Ov1N9GHYtYWkJ2TMf2Y/2zhldtYjAqYtysaU8seLTXoTWaZiA5DNSUnC3
hMrcnrOLogsTXeUHb3z/9CelWSVwDXcEgd5ddnKkSner/tYPG7TFgDBaXdoy
FWKHbmZMQFSAI5204KiCrXWmMPYl2RhCZUYbqhwlX8Hm1DgYpNWArv99E68n
Sv6k4sW7OGiNv+FP1aqMLrHBjh5asilgmKn1OFBavPN9yeGY15jKCjKA2FmK
XCegjIS4z1wRR1dqDKwS9QBhxek/42OFFgl3QH/qK1tySX6Jov5lVJkxw+rD
DLpJ1vEY+Vac1m5K09pnyLYxsRVUdAjXti3kx2CVjZqt8NjWkuxPd/RFSnGh
QPsqD4+krP+UfFkUSVaxPvltwiB6AU4y8sTyUSTwjFPMUPChTUNfONZkEFRp
oXIv+c+hSDoEfliSJjwZf4f7f5XrloRy+Us1fdABKmtq3gaPRhGlXSbnX2KT
okZesMkjRPGAW1Fn7CgD8hbMNPzujY5l25BXt++Gq8eLn3JZtffBPOn1LrOd
OMpWz/EpnPdmDP/kBFbAKeVvgPeKZndKz4KGnRzaeMhTYJjz0uq8lDAWa+AV
ht1EJzcoU1264B72rkoz0k4LBv8DmseludeyIkZOUm/oKXrHXAjg/LtQHdOY
nUBvGIs08/3/2Oc2UDuv9Z/Gk0UIke72SsxQtjyHlqnhwamI9IX6cLdGdRMo
z25lnQgRpi33ZHGHMFE2fcjv34MAzWmX5PBso0kKZoiILGIHqxlnDitazBrH
3slXmjm/TEgfcwmGvH04BR79lMAbhQtVYAIc33/uyIfTJwmGBKQOwsOL/3YX
y3LrwyUptfFMztbjDjyhe1+8kNrtl0qAvUgIH9TynVzW7TgVw7yCZgKEtZPs
aTeBZ/o1TtXDOcxy8s3Ll48Bu0zpOOvsrBbVgbLpxw8qv/PONdbdNzRmRDyF
rO4u5QDDRK6HhPxvOyhn1Mgfk55SnTY4Qz5oQlIi564Xc76hSwvs67IhEKvB
2fPUcYCJKniCw9+nFdzzt3yJTA+bRhv1Tg9sGsup/7ao9obFqrZoI6JVqo/q
F0FhQ1HlbCAhvZSVLxGYlJnrkXLA0+47Aozezry+H6AnqJOCl7yTJSG+NayG
YoB+7cd8F+nlx7/Ns8S43SAZ4DRL8d13qqJFWMy9VWVTVZjhiApJ4HqO5USz
PZhbs4KZAVcsLt+6TRd0mE2KIxEoo5nbGcmbZmKdoUxegOOi2LOfj8FmFadY
uq/eelmjFrQLITqPGNQf6JzV95FZwLdIaHpMzjY6eq+bq7M//UfWfYj8fs7v
kI24lWF5IBZ+IgLUDARxtbqD7iaIjjfWxB32tPSiwlmv3IzmUFNFxMsLBVMO
aXJ1x2i5BEU0DRJFAGaXYZn4giqnnnHvnErw+klvfPt3TwVED+E0bqM8LxR1
iYvJ94U6vfB8OTetDAPn5xYa85KNow0lPFP+VBhYDyKrbJBrLpZSh0U0JC6R
W4oVVQCQAqGX+m8w5S1akGX1Php93fXka6ugI0G1123mWUPrhyumjl2H9MUE
iMy6i5fNgrg27VMuc6JgkATAw/fOcfOvQZPuxia4B6XSxQP4O69zDmyGvdMK
EfJMU9I1PUMveXioKWJe4hsZn/BGtee8KKuqpIygSl/y1XoBbUqSmlh+ACAf
XpYM0BHK7n2LzgzYKIDMY3BuATqYNOWWNDTXnx9T2hJPZeO5DC4KbAXjYgTG
NV8vOx/W5Z1V7Yspdbqy1guwbd/q4huyX4uXIETKx8iLQCxHm20yeK8gUNJx
M9M1SnYUvPref3CF7vZWOFjhtSdwEbdtn2glj4p18tTRTMzkj9kPm2cDXOcK
P7RHJRRA2Njy+ftZ1kyOeK5sy7+csn2iE29b9yxQWCA5aDj6vfGHBATJUoTB
IplBl3i0A4CS5PNaKVwkV51enY4u2XZtbPBoG64CGC/rFXtJEOCokBziGncu
RYOpBTjpxyNxPzmIZtVfRaG/VQ7WvlDYFHT7/g0uILtH0TbFfxL0ZotL/CBc
N/93PpWPvl767mTwOOdPMipxZHmlvwERbRENeifL24nOBbEgO3eGRUabLB9S
utfYkdfaLVcFB9wXfs2KChOMFnt1nfRouHm0UXAwM9yps1QdNN5Pod3pmIQE
NHjo2lB+vA+k+d/pnTtHFobu33fAKlixd0oAFYJUN3oVymtT2oyPc9WsLUTU
FxeFZLcjew9caNWAk6xmwTmBKHMYoRZo6/hveq6+HpJ13n7cDB0UAXTo8F02
8rCpLtfqFGkOweTj4ELcUeGfy8CQB1hQlyGXJpChPqsgfgGP1tNVF3MlYAFF
mh5ftyjpX+xRinrUYP9zFK/9M2kBR7ojqum2ciyt1R1RRubP/Oeq161dT22Y
6ctZgM1RakWbmLuhAU2gPt18oKC8VXDeCDddOKjVMY42Tq2mGQzxTX3T829d
IenF/QUx3oCx8o0/ygVR+PRx5VUYMlEXATFD7YD6nQsMiGV63gv7IWqcVqmC
XNtSMz1PIt52hD0sD9Jn1/tprH7El6hrOsRbSnqbOXWBt6UN+zPmtXxcYDa4
ghICPh7fLkISUUnHvJW/35zdmkTKq8GBZs0M3tOuHvFy2xLpNFz5O9UU7gsj
mcNBb8VJnwKS0zq+QYWQQ5i2wfiG9EEfiH6YWrcbsR9pvh6Gb851nO0ooj1f
a2ypXi2N2qMqPL3N7FFymZ/8qZ03Ndqz5vnuQyJCNXAFMF32A+U41EOSEuFw
tw3Jd0B0vb0wzH0eQ4BE8e0wypj9zelaoKBkR7INMvW921ZfEhWUUKSEplj4
gwtDvRlltZ1ZXYb4qMNLUsFstIYlE9fvGS9Ka/IOP8a6fdTKGX+MLzZLZ5J3
r9DyrPhT6CNpzde05E79dVoesU2gLZ5qVhsUL2UFOMa9+9+DnwNdWiGEzcnP
+deFfK6PZmbnoksx7W/RAeh1dCThtNeEAyvREiHrfPyrjxsXrqSMy7xHgVhH
cUjXMFYJbKQRHx0qW4b0UM8daV8Q5RXpY0Cnv9czC6gvSOuUqMxLnV2DmisF
4+F2FZLaU4I1agHWZ9rLwcsDfFGOeIzy+F59lzh4z/yeaKHkb5HUl3ZNbJMn
kFnnIaNqvzE/8kTFPRwt5iTr/6W/tGtR3cuXuKWYE8PaDsnmJHMdWcMctEkV
6RwzV8TnArxnt19wzwFimoVMLHrtMoMFRkcQMCiMZqwqkkthBnj3Buf2Glqz
tcCXjoXMkgSINxfn+1pJ0uSSDk7Ue/CZVntNWA0nT332Ht19r0u9fjQVbtiR
uuxARpGj+A9cCeBT++QvRLfvRZGl8UJnjVYmAdNbUOXQxFVUPz5sgfT5pTl2
84LLtMP9GeFoXiQmIFpeWaX0jTxDXJMs4MzQTGvTm6HbJ/97pBhmtL+QaYVo
xyykXEvadkca0FZzdj+LmcWDFzH9fgr5HmdDylBcAgy3Q7wvBgF0XxfJMd/y
x9uLn53i1TVVNLCIQgOg7/uJvkFyJ3kvT8vc6rvOSYXHlLDsYNLh/slxc7Lj
9tf0AyKzjCAdjs90lDD1TXzTPD5fB2sZNDH9W77o9BOiNfmX2rDHX73waZIe
cb8zZl1Xfd2OiusxdmMfXig2Q6R5XEWG+IeF0pwjGXk6idH6spgv6709Xica
aXd48Y9rGTLT8wya0Oap54X9S3he642+0pImTU7iQQNsNJe0PpimvHHexee3
mKObENvf5SnzLKQWTwsOPz9dNgHhZLWqUrDRpfKqxirDhc4oT2jw7QpdE9Nc
mSDEp3gpNhQqExLYJ6WyTPHa3VvZuErM8kARhBhJQQNeYddjL0DtaNgK9+cM
tgTKpyi1WdacHbK0r/ysnL8ItOzJfq/kh06BHZ3mfbXqHNb4bY8bTirXdrxQ
vAdK/+j5Y700Fii6UpI16FIGpv4h4jUSXUtYOuUl4Sn+Hue4M0NVhp6CU/07
bRQJbBUgcRUMQFvLbIMBx4dDnkoK9ZuXxPYDUy8i7pryiJemUGcdiOcRQgze
X+wulDjI7M1qLy1c/QxWh+PbhL3xb7hGZemwULm5SxdGI2TfS/hoSiHp5zHe
V8vayd6rzOLY7lyxoPfJ5p3X+9BpJTy6jhlTiA8ba7olyD34iJijL3o3fgK2
8GVgjTq6KET161Lt2ZJOjFglo0T3IxnWS+vTC30zBvdayPE6yNFpI6yA5McG
2i4dkVdVG7jMDHjAU70wLQZYIqOp4Ath8HZZ4ZJ1G80uBlSwdj/obsPtX4Jj
lP8HvH8ZwmTXLJNFPmHbd3+ErSofrfA04XKfqdM4zz+EYpK5Eg2gfkU5Iebf
4mB12URGqqkp+BSUJnmPfrPtFcvlEQalWvFXqa73U+DHtfcSrRZCo4Vf/VWS
qC1hL1pWbFet5/9YksRCPoe0eRG/WrRwp5cdgJBgQxnSZovsOY2v6NYKRUem
eQtxVfISwZq7B3pqHvKHkppGNL039IiTCOBieEAIkhm6s8G4aI24aexI8HDD
HJd4nri83fnToLasSf9nfvCfc1YHufCwEE9YVxf3pZ9uZT1EuZi/i+XsjqoK
h10S3xyFwCp0/WXDmcP1a/kPfTFnEM2PG+HAUU422VcSuUJfrk9e5rQwP2zP
jy4tIihMaT5eGUZAnuiExEPsuHn9LcxBjEvk7mY8aWjchFrzv4C+WklBCWum
lfQR/qYpq+oX8dJm+MFNv/3C2h5NL8SmhsQu+zI44Pod04v+OAiHdRRgZcX2
BbXP9zAhxvk56D0pPNYXtSrTzFUR6vfz6WAg0GJ8MGjsI+idD7aWRaMsa7st
7FVvpFurcASsmclbD96LAGkzfp8T1TMubVqGALpjze79w0e+hoeZdwjhyGuk
3gCk8MBiMrg01FxEfM0HHBHGBr4rCY2jEM1J64udZAIGKkpUaYhVeP1L6Wnc
gxumtHwTOxBnRk2luEQpzGVCr5npBdeRRtV18H+S5Luf8VVIzwcx3EV361ET
UJmEFqc5XPY8KnziLRs1XPShgc6SKgZ2zAtUqGPLIjtrtPH0XrjDQWzumvBA
aVojBITpN3rmSNS5JenmsEDYuFUO3zHuKzTLLFZr4ax/aKC6RxB/0Jjuxwqh
Cv/vMdFsm0dfiZDtml18d5EUbOxYGob5rwIwPlXToLZY1iI84Dz3mpGZQ4+Q
5tdVqVVeIOCGHiVcDDpWllGh5DobNvGZoKHQMPpcF8fKsUenQyeQEbTo0/bs
2Bhc/d8cZRsJkCiNGoM1ME8Pn+RLsFwrskzSv+xMVXG8+lsm11bfqOX5negJ
M5CGzlwuELU8WKqdOIz3vahzaqSMghWnDa9dZHcTOZaKY/MAPP+MERpM0G4/
Bd30b2YwDV7S1fnAUvQrVaGQBQzrDP1wikg5ob4fObfnhjqUWJbeiw5LfUJH
NwTkLNfuOoU1Afl1ggbEY9eb5Rrkie2NkZJ7pec9b775jX4VXAkJIwGPEbxF
TZEmAQMP/qb+97lp89WBcEbwBRPwZAw3zpbU1hKVK5g8cUUvF9Xs85g6nJDg
RI74wFZSk27BmtvTRP9fDPsKs0S4X2ml1cUuHMyN130jtxlmtARwwQZs7HJa
FYljyDny60+vUdu3Gyd2BB/F9gv5Cwf4XPv83U8RaTlCzmXnbE5SeTXte94o
3EL1cnNfBsjSab+w4sQjfQgbp1NmtyHVzVUF/9hVyJoE2Vhz0LAMDu5wJ0TS
hXKIVPKLp2PYWMb6CI8ThSyWqkNaEQmuqbNDQ6ONnXBQj06v+Q82wrvpiXah
IOcn8eIuPr6lLqHyWMK9WUWntvYRJGIC2WCT5mAybfovvUQXEYaiwcsE1nsy
5PeY6knoDFWlro5u7YknbKjyvwH7zd3el0bPHW9La6A6/YbHiKwLeiYm1OdR
ZVgsCgQ8NEgsj22uv/qsdCu0fdByXm+XBujpcph+p64X//tIODeCSwoWu0qC
2CucSZ+ogGfNVmkPJaaKnADnIOgBPVOOtLfQAWoSi/gkuIfDKCXcAvoNje+A
ZloDQksJ7tjWH4nuIkoKbagVeOjwWTfoVtcQgTAF6rEk9lA694hpX1bpiXRz
vxBbVub+A/gWjKfUnhnjF1W+e8JNVrWNy/4EVvy1SnXK7bBBD5XR16s4vsrR
7ZIHydb2+ee6ywaWHxAEepOGnvsCYk4bcYg5w6EyCDZdnDB9bMw1nwQxv0Zz
8VbsHT28KwTm1nUnq4Uyq8c7e8Q9kgVW2Py+z1KHjpLVmkz1c+48KoRWag3A
wASy48G5VNIrJr/V7BF2Jf5eI+z7LE98TPkYiybCm1VH3L25tUYFi0E1EEit
g90MCOFnQwNB0LZoFUiEsP6uWoCsjK3S/0ckjq4QdzoR5xyv9+CefGV8dckE
btZ3twMp8W6tnZ8zOe6zGXxf5zbQeN6awR9JUrs+lF5WdeG4INh0gUMn/MaW
d1cfCbF3viY2oePXDl3fclDUyO0OS1skLFRm+nuRYziyjECg93+BAqE1yMCe
gy6Z4zYXTcz2JGCFfBdofUlcTyHy0uwbCaigQfXJoSxd1Qun0OsFvyXdAquH
ZqT5LoJFwH2P2McZVB//gjxX3SxJH2wsBaRw8+xs66aoOEI+7eeg+fMAH6Y4
eSNDcmof8GORHQoD6R2/Z61wh8Pq/1qRbXhdHUPG/l7dflSmiU5JCia26HrV
O58uKX13OnYUXWq53Xm1k9JZno192KcqO7e3B1FF4GMKKb5XmdmHNHAIb3AP
PpvnkCtbnLYwK2jRq1zKN46Ks2schZX6znr+FkaNHoxP0r0VFbwA7r/hO1Lk
R+XDegz1xCQiJDP2pyhmZkAUHiNec7IbdnMY7YpZOIf29Pnr4EOW9LqixqPG
/M56mvp9ckxAuyutFasjXX3MGcHuYDWDyMhnUKt6BPBt3S0HcoKu+414Ca9p
GgSA3zwP4wRZhQBxr2R9ac8qhMipWD/Iwyy+DqwkVIu+Fu0qNY7svgooprQV
v2FMU4nNFNxM/Pxy6nkiU13DIzhd3I5LTEhYZJ8vekgLp4GxM//+zWwk80tG
d4gi3TVXgY4E5AMf3GCxcNGxld/syzyygOPrLPXPHa4C3fSgTeMFgsnkMJvq
ch9GmFyW3JgMNo2Oov4bDJ/WVI7+X47NXIdpjAiZX+8dF98p7Qk36zSwO1jI
UvH+QNEOP+/lMEWAQ0fflB/CdQa7/f+0zVpPTLvb/UpxKhkaorshkFeA9XOv
l3UWXWq944v7QpZ8um7lGNQx80soPPO6AtReYFM40kH3k4TEqdT1QHF86R06
4fWsDptUnc8P+r8OZ4Xdy/w5cvs671ngnwhWxcxKCGzP5u2DKwuTIxUjAKYq
nwZTQ+kE7hjtgRN7MHOHAd3NV4TPEKK+52hy7TX776yZOFtxAR2seCWRZl56
Vs9oTxuIbKg40r4zrRA6Ku0FDouO6Jc0Lms/PVMQbkcobHDygnMJdvCu+MPF
d6X1VWV7sF/4Ab28rPkBB36qF/s/vJN6lNrPKzRGW05fTj3kKGfdF8BwQMxM
bTNgXRcGCldDlw3kYSRrx+iM7TOAnLJxDXhXTeSkPqM9UFHei7mAF+2xXbSu
aaKNcGj6QptAalfee0pFf/N+UvJmgsIt+4qJZDiiP2xUztrDamMwakHKvG30
xUvDiVyX+3PejfZS7rtuomy0U7Efhw6Kik2+n7NueW7sFcaQzVKLpDukediK
8MXyRV/NT9amwQ3d38QGnwfnQG6VXIdg6JP7wvcUJCuXEN93BEys0v8KBpDm
ILAAtk1DCTTjFNLt65WrYPRWM3jsCadp7YyTgoH/jhtIWo16a5NPxktz4Zez
DH26p/v55QS14DKjo6NpvdhSyYbkBMJWSH0+Uz41h54H9/Yfiygbi3UWeXvM
PPMAcqbNWcNVdWRspbC+wyClbNb+8szDGgP3Xdl71I0crPjLrhaFsEROndy4
xMUdusJ4kUgeTQ/uOnrAdhrxDSZPe0dhPji01HIwQuJpbvN3OG2txPHMkVHA
XH/icfN/CHmhi8WD04X/3bOJz3QpuClvZF+MlvozQLZjxWznBwbascemWQqc
N+eDlikIc8EJ6z9N+RMnxmDeyvNOEA3ltyWqZPuENvTsQSGcmCmdO5vmZv45
JDBssDTGtmn+djGdIg8N62g9sPYBtAbK/DmLY7/9AuJd1JrQu0xvMoXzq84L
65N/UeTbHWTfN9WDKLVqk79ouOPQbNWAFInpRxZUXTXoltzvUB5KMRSVhwML
ttYLal3Ne1J6eZUHHBX4LV7dsojRMB8z8Aa3+1fRr6RvgbGKduY1i72aRAg1
Pk/H6sWxJxOpoiyms/+NpZfEXtT83jUgdz/nn0e9+9yxO5n1vGLv+VrAZKAq
ywfyJuEJprNxZZrcR9tqch/otTrwQ5Dnw538rXmR1hWHEa8lwQZC5ykyjsUe
aTKAkYbxJOXpB2HA9LW6XKfh9zoYSFehld3qWeWUlx7AFQtk3ml1nSiqzISU
3ocJqb/L3AnWPXPemg0GGJUAf+Xgcl+fvMPrrW1ItDBOrc1b9WqP95Shzh53
nfpjgcLf2jZ3KbLH/g4Q/bH5f9NbXsMEuVTlTheEcaC1UkcBek97BY9f5QnC
imdkhRuDHsHH5n2OnbFIzlbb25st21+z/Tg/b6+SeKWqA0waGn44o5phML00
NEDfxNBrhaO/eustRKRl58nk4dqWyz8GnxW49YCx+4gYerCAsBo4OKET+T9F
C09L0ig1K0r7eZyxPyq6j69Q8YEsby0ncVTN/NgDQWNTemFNKbJ6gUbOSihQ
0ubtlKF/DfFTPid40spCeIFoSKkBKli3s8xQLqQ1/kfoAXI0WBNChVdqYx7s
acqfkgWjX9ql9nEuj52K1jutk8+L7OinCMvyoVRADZW4RrmcZ9KewtDRGNZt
gOTScpgTUYHaBm3f1dFPhScnDT22edYONeeer0pbTiFygyQ00fHyJCloGd5t
5YDKWgWZfkFOMCfvyPiV0ISwHfYepeaz8jv0UbFy/PKaZ0+ff1b+Xw/l42VK
Y2hd99roFO968NDmM9Fj6RMAAlhFOXxB5OpCzQdCuZZRdzChsS7QKLB+5PEE
OqmpYmYBcuZpuQT3FMWO8Va0FpOUKI5qhYVzmTVw+RNEGvu6wDyN/hGKmJ1b
XtW9jwNOqj/DxdDefSID8+nEueZwelFFK3J0kJRGpL0+a0r+DqPG3FH5waCm
hdLi+AvKzWcF19nCo3gD4xKAnH8eJP/3Gx0tmngwnCNI45Vp38TbDCAdBngO
4YgAdUFdO/uij5wKca1RXh4PmTXcWK/vbSicZC8dscG8Y3gg3nRjjAZfHBgC
T80az2dFOeVq4JX/kuIX50AwaKBDsUCPgcSsqMm5IdsP4CrNUW9RdotO8yQe
w5esn1OwbG533JCno/xk3aa4HH7jv7xneo58Bmbdz+zlvv/tV6cfxSnWp2Ax
P6hDP/8JAXPNJJRjNmvSToqT/meQBC4JdZI/wWPUyWx7RD3g6dfwi1M3fx3N
m1EgpSOnqT7mzCD6cMSa555ymgl44QN7835yFLS5j1/c9//c69Vg7rYmscJu
0dEh6EyE92Vmb2snOFzMSiOTjigp3WlUz7SbLmts9g3yZoE+9+d6l6Lfm25q
00PU8008YF7Xl9lvKS5SgTnXFETQ1YTWyLEYzR75thImQoZI1rO9DXN+9XU2
+LjNclGh4WBXW7vgE+sR+pIEP4FPw3by00M4wP/dWsoB0v3QF+Rsfm3pgNpl
17Ad3mtFJTM8EI/DKqpdG7XhpI2MZGhUmZg2dz+hcDajJbf0+4hukOvyvbau
VmAm7Kbfc0xHpyv7YcpiwSHniR3JaSQ80hn1vVj3dafHNNg1I6dnlLju+htK
3yn7sJeedItuoQho1nhbsRA9Mc677lSxNSab033xutPzgRqiBDidm1mPoG3Z
wf3NHvTMlJYFHE+YG3CHVbZPkolCrZTCTS407E5fQO5fIseZ0GL5shTltICQ
jWS4E8xY+jyjDMgA41uE5e+jKQG5vvt6vaYROobyYEsdnfkbY18bzGoYGdoW
CtjQxiVJ0v8q8hDNfCOKQ44J37kwaSfXaVL51vEhH86auv0+VyYpRC2Ncx9U
QMenJWvsQeJB+00n62CHVj235MohXTbDg3pCQo/EYPMgNuyuHLVNgZZNz54e
1o6d/f8mct7UhGKs/93WjVl/jAiCOn62UdKB0XX/CadWhkYTXRjfza6i5EeF
Rbepg3lXLJCIjh33cjmERvsp/IG7tqmQ6z0cC6ZK4yQmSFEPLOIV+5GxJ0ct
shXgdKmwjsmL5bC8O0TfY4HzrrwCTMPRkBHO90GlYe7yXZL0Apindfw06hvV
lYIwo0SuskOIQz9h3SME2MCX53lC+r8MLcDnAtdjnBdv9mfGiH6blNwvNZbu
rpWr8jOMzvkdc0iN/XBr2HCxWdnQ+9UUMwd0Le0UYrURTPTbMW0z1G33WfTf
JgjlwamH/HYtKMOARQREBC55eVCZPVoZdw1mIFYPMpFdnoYvguQ907lkSI1F
TU/n5GQFnQUfiddRZmvnyQyZRU7xdHWA484RMbDs57VbcwoV9kixVC4c9zUE
ct7IEnIVpBvL95B7rkE4urKSBsETebIN4Oa/qUZuZYAmqL8PBwfMvgo26A90
lEQwjtcY82Wuh/LLbZuhdO+ZiKqwSJmSPWuy4nIPjifcf3YgGXD30byL8rnd
EJ5JtTHBMG+cbiwtmQhrr+5Nra0znmu4BNS1FNskFaNBtG7ea9cFJH4i26iY
8gKfoLe6AXOVN5Z+i3AACVV+7E05ujYCyhPZeqdPgmbYy/iaJkFS/Fw3q11+
ShSV58ngm5sQi0AeAUHT1iUGFSc/p3FVuu3owLiLLZcU769VE6uBG6Tavyhd
2wri9xSphbGkEYSoK1eaJNF4St9TJK0G86V8hWfd+puQnNXYDIU35PCL/H/k
G43pB4zrB7VOIBrk6anhQZpt9+pEa7zV/2FcKYqmTojmkGEf7xAzIkN1hS/z
YvyMoqhz16gt5f/+Xp1zBq2H/8b0MPb760FMd+OyKZqYH3gg+CYL2EM1rdjA
gpdGO0WGFsG7KQ8ct1iIs02PaeFJluEDCNo4fh2cVkxavfezcPLW9v5BbgMG
oo631Kvt3OcJBH8eCGWKhKUiLIxL48mJps4DHLma40U9bM0NjJpJQyLK/qk2
rmkdrIiFMc6bUYQO6cxf/qyoNgQxeEzNDnW9EOUfIfO1x10dRFozYRQFS2NE
fMuTIRiSlaYu+TEdoMpJcKHyyStjTcubkrHRzSnk2HGf+wSvLnFS7qBRy3/Z
W8aAxB5YCH8aZvg846mdgDmgT/9BXXT8VDbKFdoWoVRS2wQ5t9qXT6Sz6n7b
IY1v4jqi7BzGylJn0z1ksBl6yZR0LIkXBTQv9L5YTra8cxy+23WeD0+LLGM9
FZ2c8S1+QC2P4lvkrDwkaXNmEbuT5VOyVJvBCmNfwp0C7e49QuxBgJJ2IxlO
AqVEVm72rWYaxwEisbGQrfnhKyn+GWYZx32xRXwkxJEy7gHt1MX88S1XV4Vy
8lSNzju2zVJlrBYPE7oGr9yj1AIPinrXYAETLteigIa/TlKEN/yO8HBvtQRc
WkWiAtnTk5CJxfCKGNvIo6AcPb84a9RGlK2lDNLAvT8HqBQLy5x2g3r3CTx2
CfxFrOk1Z9BANvnXJKexvDalGa9wNu7ZZM2oqIeTVeF4xog6e9WiuDkx32Fs
+W+x7PBpe538T10Lxh9AmILrzynEr+uaR0HEFGloRj/PGZ1aDt6RkotE0m2L
+d3yJA7lvxW+Ij/6kKl+ltDIp9neAYW+1iX+R8t2ZXRYOQt5acC+n5OdOJxU
LmQinaS7v1cNo59ZAhPP7bmtZYSA3yajfmkdicCaJJUcNbZfqiKbBAQ+quU4
IZBcBFjvTgA6bnPHvbkv+d7PnTZlSNZAROOf7ostt89QT1vNIb3YsOCWogdm
kzQqLt+vERZQuKu4nybUs9Fzx10VGj4J433q2lL8BpDBZk6a9xmhNP1rRCbF
Ursii7Wly6rTloKvDIG6TGcADSEwwuXJ9TvbHHjSLJSw4kI2IkHEfl6VBOPN
IxHS0oFwjWnrfT7P3z4oGxweLsaEd3kpNaF9u+paavLIn/YYEzVo0mByhkuq
sez3+npZCG9eu/nJp2DFoxKfrfwyN7tu9bjIbTqEjyZAxrygBGcZ1ZfPlaKD
VJsEaNToADegCaklUj3MDtqmnerzhkIwolViUO+qWGIwSX/Muy+hkS8g/Hy4
nwn1vk9wwBhgd6WahnonO6dBCCgTvQGovvJIjHgPSosB29proRrMohFiVifX
PZVyuM8L6QUyK5oBo1TLsucYFaMoImRYLkGEzjK4h3yF5pVDEvEDH+/6aZd5
J6nrl09DDCjlr4lTn8zeEZWDhKSyLTj+/oEZPmID0E5Z0A/3DThX5p6aT0TR
OKTpvpF4oSmFif2ZM04FT+qFPi9zdxrtcCEs1vmqFjEJ+ro0BtDDCmFikccb
C0fD/H+PNOZNdj2ZyT4ZVYQPB5JDx5avOy8edhf8rGJG//xx7kT5uYSGkAyy
o6e6bdnU58B/abHSRJK36ziFiG5X/FoVMwKHa2PrttYrCs3CO8xr9hWXVzGF
zkjMDSuWogi139sasySJM09n573YMR7hiQ7rBasUO3BYRip+mHE4YXsloyha
RvFiXy9QC/Iw1EpDJN052vr85RV+3Kb7zX9HNUz61InyXIZxunISslaDdVpf
qJ78qzAhqca364UE82w9AP8b2Mccoxxhwu/4gnYkE5CNc/mJRVztCM9qgglH
tWS0Fk+1sIo2VmvcKuN2f0cu6cr2OeE6HDFi+8uR5MK+ZB/cd8oiopvyfbh9
2X+hDUkeYXqh4c2FIz5ypMoXmTIVIIMs3hO19RUb3IvPIGd/+6g1QgpEwd4R
EioePzu0WlrWmp2y22qi/d+QZLmZUDYsX8zjmjIkdBEvhg89YixmeHSZHTHY
IeaDv/g1rJ1X47MRJP2FeUvLshzUd+iAErJEzvjWCbcyWpYUHMSnhJ0dzhyw
vfqzZOkErBnOrZ6tyNvGgy9Li8Zl7pH3yz9LuJ6WfEsB6mFq9GFpfWbBBb1C
TUpYruILFzBZO/SKAygh1B6snVH+srr//rD9lY3bI4hlYesF23RIq5b0CPQ2
KF36D3MLHbTTS5XNMxQ7Q/L/H7NGhOhWhbnfT6zeBpshmFJiM9zm6seOFQMw
oSNUF0OvwAQguUTcOHGA5zj8wOsWeSchKeGaZvlblNiesppuAuny4A86SsAy
6CI4l3XMyTR38eyJz+UtSUtsJCCToPSPFGOsrxI+XUH+VcJjJH0J2PdgdtNI
BHRaOgX/WR3S52ayzdMBrSdxuSHRfsEjovdmkAeY65As3OmbM33fYldn+KfN
WigdO5IryvoL0JLl0OlCyir/7sOoRoNPmFb9Bqh8nV0B8Iks+myQX8IAOlnd
EpJ3CR0jPLGFK4v2JkdVKYUdntdNpf0jE6lG5oi2eNUJc7UBKvqYPsDSHR4y
a+dNA9eYKC/TYKS0tZWaJ6Kf3CnJ2yKPrxmQELzOONNWbvARQkXelKteztbs
yDSlDzsTZjI80YYxZGKReXwp/K7QAEGmnsUfhz+fCXaK3C8PrBf3QFNiG54l
/kYK19E/S/d+Jm341nDrzy5rSzl6frOSo8bAHAogjn2sPMw2+I+aPHti9yA1
tGoqh1dZaa88S0DxrYD27XGPI6i3IoR/lqrIGF2di/OYR9QLkHmGvHWvbvIh
6SRF8NPScYWvtUmdIQqKKESHAJX5SPcFx0hQRH4+iMFPMyJosmFUIlDFH9Uc
JvVTLtVJ+GTeX0kOo2kvu9m5YQRCG6JV130jQ7Mda1or5fEMWPymGtTl2dEX
zHJI0lxF9R+DJZdxC5/K7nnn1lKsCfBNwwastptMkuJV9JlhgmUoB5zpOCVS
KLSViLbISJAyq3SleQcSrY00DoRWPr3SNsWpjGO3jNSWkvC0qZmdFT3T8iY3
malZoqk3JVdgz8LRksa+bc1+8Fqf2CHYToZxFxva+ncMpqHk2F4o/9CM3MrH
qgfqCcoS4xIQqXl04QdixoAKxSNTdJp7bD3l4YtL8IDqNW2QUDRBXDPP00Ot
ifIvCFnJPuKE7KGaelJz8gV8N497Z7wubmt80p8ko2JnZOGIo6QK231n0fEk
Nrhr4tpyIQ+ZLA4eagbff8zMq832f8/cYe71imhaugqqXiZsER8KEeYROTya
sTFB3rqCL4XEZ7Y2tMQfQA0MCpp8L/s+WiZE5RcSvpqxQpp26bEtWD1ZkbnO
5YKPENrjoy+1ZHEYr4TFMa75MIohsOaFGNMuGqxzd3L2xwErFlAqZYGuVLCx
Z62pndplmCZPqbfCloIyLCG2PI7lIpc+kl+t/eQ8j4AFfVdhXW0hYjuWqQ6E
raXlYDO76iInK4KpkXTXBWTkDqO1hDawqWVSzUmwjzuTh2uG0EffIF4Ljglj
5bMR7kxeIQt66KEiG1d1jgA48uKHb4uq5OKebg5fjj2NNtKvDM2xu0yiwZKp
UaQ1ocxkY3mNExy6soZoY3C7HSksfWGSM6w2o8YBfLfc92dadZtkWJsoS1k4
jdgsZ1yJkRMEjLyoHsd+KzSdBrRdqZ49m9RJe6ODxIgP4gmMANvGB2Ybl3H/
h2LOh8vUs7XhcFxCAAKlNRZ0IRr6g4oQmswpN/oO9D/LvxUyao78gQwN9WEu
0qERLl7/agPVDSoZCAorrNFn0MR3c4mmjjsCpq7hVSCVj3g5pGWNAIdhvYSW
7cqqSfxY++I39vTJOId187/UbDDh9hJlqrbkcEWkyg/4XDAH8zDr2qApYLQP
991wd8M/ia3WcAM1pcvnEAFCFQzeRKioy+Zjip/DqThpDdg+3cfA63ymIuax
We4AF+CM8nxzpXQDpWPFk+GdUqqTg+MKj1z6pfBcrQLl0kRT3dZ6uqt7dhvW
LF+Zx2CzLNcwRhZWzVNa0Ol9l4B66ucH27E/ISOGvBaFFIG4bt243lXgonse
03hyvt9aEX8QmkFyHe4NjinzaOE8QMA75UvsTd3jNhWHYUPZeySRBiEAAD98
QpkdYkiCG8vHR+9HPXDIGY8OmjZIFwRXCsg5Vf75cB/QAw2RRqre3fDEcsTp
f+T65MJzwbcu7qCACSW5mG7kctkph79JAJdqIacrsB7VgKFMKyYVVDw+Z789
GT0cfrz/cSP47OszGxWETacuPItpSx2PYNCBZZP9+Aue6E0uqjjQqSq1ik5e
WRLjYMJGrxsMKBS7s53Ign8oEjHvZyuyhiOO6NUT0b9SexU/D9g3AV0NNup0
YCBx7z6NZjOU+aVkGF/WERW1AtvROFJun76MgDmeswYH52bm8Jyh2RGh3RJL
oenC/pa3En6rCEOT++oleZJVgdxNiRb5qvP5/oVTZvik5aQaIocK4owm7acF
u2IIkJtcUV1bZH4zn24EVJonzV6oMv6gcqJGRxHQ2xgZixnLaDoq6/YKD5cu
ZaEnScb5JMOZsVk0Et5ufUtWMsOqUQj7G6CH7Tn4yIPxQJ8HMs10m3Sk9rCV
PBLQ9z8BAztwkDKPzhO6jB6cpIWzEjD1343zbryj8VZRF3VPod7ysfs0LKTr
x93JKA2gr1Fgc8f8i/rQZcZf5MvjXaLEz/PrrpC8EpO/lAtypD1MQb6pYUFZ
EQbmkRffYqZ9kMFRaUUikHByj/s61iRFQr3KtAoXuICNtYsMmLRIVOBtukSa
rQpYuGFLEcunpMg0QzQ1Ln9GWRHzy8yllrkWTHuczdzgiFpHm3AtGfPpseha
qUiRykTk0jYQ1OGHd17WX2vsZpe1vHrYIucyE5ax+dBvWn5HkJUgQFGtciF4
ZRK98VTAnl5oQJYsHL5I1rI6TlvxIsbdIR4kwkM/FdK2d9fWo334dEum9qke
dqkYw0dc0QEq9EeSitltPUEJPxb2/wZEl3vXPlLhGFjbpOPcBJg8jCyRPjS0
mlJWGZNXId77HdHAr/jWF/BKYcEw74LOxd6/0dHTkhrm/Rbu+1DoU0rvMkad
4DYsB2cAeqsBm/zoCFkAV/m9XRFSIZAAehQ8BQAHfP7/BGMJ35iYeG6qDb3Q
kqxlbXVNe5c8GfaNwNKJsFBI/O5gecoUSND5WX90jx5Ko2BlxPc65Lvwc7ve
Ctgzpy/bd6zLbRFw/WC+g8I1FBJva1/bw5LRzPniB3cpAibv19R7zW5M8GBZ
nSQAKlTZJdd0zO+JxRbI/+Pd6xnpoYu6wj+23P9pW9P9DNrd0mLGxLc4Nt+l
FcKprsmSf/bdD+VENbDoyUsz66+VuTmX8go3A6b9M4ONWtB1uo0pWXpGMHBS
JWGbGEE4dh1hTGicj9La0KjBPTfkx/UjtkHWmbADS6ACarjY8T7MIzuAr/oF
hEGcD4yYEOubnWPxVsVWQXDSUy8TYSfxhEgHbeBxyeYixK1l/a2gjIiwH29t
SYJZsHlrw6Y3Aadljrg9hsW/2WZ7pJEdFri3YojhF3Bbx9jgsyfklzDBaBVG
H5id4ekw0jwYcBooG34vs/NCJ5wB9pD51y0kMRJAk64NzKPamdNPhpm+Vrgr
Pa4nE8OaTHc7Ofn2Um/S14qh8NWDKiQDMr8hb9xHZenly6jHTgPN3xu8QUbr
zKtA/t4ag11tnvsC49650uStEx2LvqGQbW4gtknu2pPcieHdyf1Hf+23/+Li
C63FO+PB+ZJeOMitEAoHi9LbHbsvuMm4s4VzHb/H9APjKRz21GZO7HdBhZzA
bOeGwn2d6178HMs/0ZKW5HWzAaCkv2/DbO4i9mxxXfCJM87NG/pVwi3rJzoC
ZkuIwOivdO9jJqXF8wN4ZGVSj3VuftrLwD8lV6qd2HpXNgruTVQWRLnByjAb
B00bsv30Szyl/uVazXdh2fhcp41oXRAva6/Z5sY6abGZ1LABBi6QNT1udRuh
bHHYeCUN/pHg4r0izpIw1Ys5r8gEcxVhVFVU4NbJM3NLTOq6d38kc0fsKzJK
9edmpZ98+TqHClOPwHhm7zvGqfygvepfUWOpfAaDvDRZKcY5dsimJm8v00Ls
bngYCTpfD1WDSbB1INjRUwFqFxgyARC/gJnqfm8uGCPh5Y228x/x0etEPwsW
EvWcXSmdvLP5355QXfwlB7AaqOMukXqn+T0Ws6cVuN94Hu46NWqtJ6vR8NuW
T923Gh5A1nsU/CRd/IAgii1eyYx4sl+8mlALHFirDz3Q0xMyk2ymYoB6Gx4u
FLS09+wt8mYXwOGqmkM7gpd0UrPCqJXn4d1EXJIEMGIZCLY8OVWN3zBmBGuZ
ZBoJZ9oQOlzGxaqeOA7Z7u4HsCBpnAz3pdRJrPLZxfWZUJt+nKOcZJYbL5iT
8J2nctbedAy57mlkqzAl10PpDfzsDar0tKrQiRssyxo7+91wQrtfNy7MTpCn
6+vHfELOjWhiBlB4qj5KdOADM99D6PRfWH0DzizQtUJOZTjEiAoV3U1DkEEC
3VlEcZbcqu0YRH4BURaNxuKjqqwKw77V7lRy3uK4SP3kl4r8oBLQQFLcorDR
Tyq/cP4o1WW7Zd/+vbtyIei5qHZq4PQS62DPWh57LSWcbJqQJkgOtafI+B/X
HDEiJ4vXmsOA0MgXOe0vC+tRGe01vWyZMKJTJMUjl1wBK8mkNHlpifeJiYyw
vAlwGCcAS/QjYd1TVzJGY/pRE+9nK057ZvXUD7+Cc+5IxYQI1XcY/z+h1iL1
gvKHOWLvsHnVOHsCP8xGJhfPSdJemd+tHQ6g/RsPP+ut2cyCcqSMt839ZFV0
Hc1OcztdigJrtME831MMItweYGC5lZ3/WOsaw32DO1rnsMuQR3CaZlEucTPj
WItZpA9IM0nMlNgGxGplsRmnp62lin5UALRLdT37wxNauv4TvJunRNh+GRzb
56LU+Ytlhfnt8iIIKckvdWhjqikXovUxnICmHlL1KI+XNswduypBWiB8Hm6D
A/zwmwCJbUO68370NZquDACw1LMNVR21tW98SEz25MwsnDdRoUgQSzaXXBlf
g+hJNicg7tERu8HG+QFsPqZvGGf/iCFZ2hxp/AdUHQO32TSVEc3kHEV6z7eu
Z8xQo5HMTCpP/r7CuIigKeqSOR/B7cfG1Y8hKFeiWm2ptfheKo4UnLCxnKKn
bH7vVQY3da7sYkjKe+vRkO4BOJIYQwSzUNRT9zy4ppkDFsHcccAX6K4t6Woe
fIc0nYybVnjSl/ZFSL6tlwgyMqRfsdNOk7K6tcReK0vq/BKfyUe/ztCewOwG
wQS6Q2nv76/LoHoBXSd/MHVzFPm/JD7FyZ2N+ac6BoBLDoGldndpA1DSGHxs
xkCzHAx9GTph8ox3vtJz3gGm9+LNTu87xJEzSlYOmVtVsHrSwEu6uyCWV/Wu
Q+SLZvY79Ed6nI42L91xtxLqAOmHbcocO/Gm+R3ZZxD9UPKo5YgeigCvaHvK
e1UB9FbwTf8ffYnWsb7MmK6QIcUdN3XKNEQECMEP5esZFzBFx3kvmn6/FMJ6
FR8BCGHFPULC4fPDZYct7hrvTv14XF9Y5vseJ3t6yaVH0ZTtMCFIS7dul6zH
eiRL/uXiixdUdo15TqCbz9dwhXuVAUSOf4OxyDbDg26AzMF9UnEJaGaYa+Fc
C560ajVwu51fk5oKiuv4MHLO7kMpZmDhcQv+rriETXmhWb5u2PEnWw5PEk1/
EY32ESZv4P9ti/umddrVyL08MulYoPDvYEY+QjfkONXMXzOxe7NNf6IKG8nK
/W8NeFjnWR4oWkwgPM21X0+ZqqFqsIR7pYwtL/WjTssu40CM0ZMWesGmEZ3y
Sqc7NVpyLAWRVHHIkoiOQmgXtnqVLOrA2LxfyfwQvJY8GBYFhJaQML58irZ4
8DWaL69JmAKNu/X92AUKXDNIolcGc0IRVYPUn9LPD/tpdDue9+ZptbCktx7G
1uxNjOYJ6+035O40AG/B67w6dhukziTryTkMHX24CRgWIsuKuu2/aEh1taS7
cTZRGgYycX4CPDetlk9HKkpEnFsGwFraQ+1j52mxqrncMKuKoePb4PiLfzIt
PO4jb6yGDWS/GD3V6sKVxMxVgUnWbOHfZ3xIpH2s87pV9THZtBqxiS0lS3S+
0YYQbUcDQktPK/TVBYWHcjDl2/26montCI/nZI5jBTUC8xADJ8jotxAyPBAk
J2ZTxE0MqdIupFvJOLfJK7EPe7BP+MOXcZ4WKxA8xw3/7QiFABfXuIJDXKGb
Do/1UR3XtugcJGngR0k9VmBkBoYU6FPpSmNwpPyzyRohJUt/GE2mFRmyL6ae
60HW1BjCkwxRYOVrB8B6hs0222L96W+HYvOLJBwyLOCt69B2PwKSIcmYLlUK
YgRFdLfA6bXrHg/2cd7ayc3WpjyfZVSeWCoS756lRznruwlKRcQC+F6ps/K2
QWH9IDEAGR6uzv1IHHuwG1jJMkOWmRwVV/w/A5uZKEPeQnChLPWN37mFctOE
5oVBPrFS1q0tTeCHl7dNSmpPlpHsWwjkBQhNCZpREailUF2mIZLY+c5Shr0z
XTiifi7NmHlYk+pRgDZtdFgTniHhsgqMv3cjIg72bcTBnGy+O0hnZIzqimN8
jtPmXOJt+Y7O3bi1p9Wo34DmxF1+KyLZ3lfZWpNeV071ouDRd0mVSQAEjByD
uUvEwptmRwogWDWxCwZr6Y8yljwg2YPI2urPyEt8WGCopZXiaENChaux276Q
oM0kk1P7VmgrmfUXlsxQRhhjMADYM/Sx/ByNal3FDl68Efcv/5ZTmVwBlDM2
40Z/RVRwW8i/qebcBODguEopeBwGjR7CN82jgN/WrqPSV5MTMT/+gP1jH8fZ
TDldRn9TZqzN/lMsSIOujWLbfNA4yZXJc7T9Qy1oBcZEUoj4bQJT1dqii9uq
GqVAYuG+M58anxhdqmzz+u5i2V1te2UUzMoQxCR/AJxj1CcmBgmsln84RONV
Ml2rVnf6Co0WrmdWm2Dzsvg3/40qW+pfRMbFx5CU/CYXPbiUb/C34I+g/PIB
V1QQiKgZuq5KHT6ElVONh1XEMIaHOf2dpA4jYEbufkDkTqCZj2JCpHHBcwR1
wv3xSKO5enRo+2w8BpSvZPC+eaxAVFBjYAmhqVglZIaRPMFJl1JJP4ITQM0Z
3U6cIKP9OiVrvmx0oWEcOLSP9gygNfnKwCDZomtQEuaYFUao5v66AD8V27Gt
yJJZwEDnj93QnAMh37zFWj5ObXy5bCLF1MVY26wPfHiIgKLPPt8My/uW8qSO
h0MSsL/UqijxaZ/cJBd3p+vnZCCAF7eqPozsOH/4JVGY2CjDPt+hxenBuRVM
JM/cI6qptahHttVBiCjv87cezY1QzL+T22ghq8JHkNzSIy5yFbLkHsGjJAWo
GaQPEEXcBDzkLnBb4neb208OzjrNB/KCKCqGeq3cU/LYqzE5W6Di2QGAassi
qBE5deiCiMFNAac3apTk1dDitHaXdftwZsI3kPov5Q4Xd4R4rP8GhNrGORke
OZeRY/q8c+f+wjwioWK7oT3GZRGfCLpBMc3EH8l1lsjvLXajrPPXijXX5L/7
1kCHLPL5YypN7xbKR3XNg0rP6sRKQW/lqiS4VzGrdnJG5R9Uu5t7D2VTyXm7
h87vA6Sl0YIseRdbp9tuiowWRr0NgKWjtHA7FoYQB7yCLvFe9Wdis0rTBkms
MeBKr8QGkce8Kw8/PBAOgVQowOX6V6xhIOqhKqRcdd6ZRWIXxUMIuK3Sc1Ok
eC3pcCcatKn6wIb+zkEQJ8cFK6rA4OqK2Km3n1JToXkBYc/X8ZGLNwg9sdmP
PfsGT5AoNh25u240xtxb7ZarXjXtadybnUPkoYom9IOIKuNc/OxFJpHvrnVh
q3oijYF9g00mSabZhD+QO1+S4jVGdNSSw7rXcLTJ7xW/XrID1z97o1nWEtOS
PSLDyCnoNp5LD7S/mBYAgemK1GSLoJ32zncuG2qawpFNCAOTo9om8FCaPS5F
xIN8Gvy/t2h/uhVuoa0A68l7xPNbcohGuUb4/qy1nFmNPLCOaQuD+UErp1aK
j2ZsZGOELbZ/2P1V2BaxA+BEGHwC/IpS7G+7Ba8mxjEfalr3Fw+QiGwpld8f
hllS8TG6vUUWhbRcrX0LwNbodfaKAOyje+ONjruRTXf4m1z7OMY9BaaquvWr
Mp5oBsQ9rO9Kp/rUL4Hn0XwyMtwWEKI6iVtxAFPMPlI5TTVkb8trinPiEdCW
ZtMOl62JR9Nw8vFGm0pjmqhEMcB599h779sdtGT76r0buOkV3PO2TTIgmDVR
KYRiYuZXGWSFt+M1mKy/MLXGcM60giCS36LoEviFLb6b7Ukm9yd1dlaZ1DxQ
PIJfE9p3wQo5mK4ZKduRLw7MzMGdyVNZedlgtgrR8xBkP13VkRfTbNm1gwZi
hWBy5q1F6BY2ubqfkKeJriOfOCA4HzgO4caCQQGT/l60NkZaFBSNt1Osnyep
3WQcGPG8puDJWaciqJ6EsDp1hskD4WFDh3XXC6udRICIdoczkkCjRfNsc7to
2Tyijdytg/pNFJtuHxyUQp3CvCsojzMPQR3WYTTHi7FE5tLH+JXgUojaqPGt
Hsg1koUUyN6ncTvSX6NHE+dIbvN0AxAkIUowsD5uiJGvhL/xUZSU0wW5rTy8
cch2as7C2cv2stJLtTB6M3R1ja0Ib0q5AKRXEp2M1MC2w6XsxkfBmwkwsEVD
Fm/NADN424fY8iBCZJOeVKC/J8SqE69MbZ8Hc/HSmESK331Ww3rjJ4tQJM9z
1LjW7iL0HN1UMJshAIt8I8p5vmo9qQNRJUnmpbWI7gWVNbIlI6pVQNuBuw5U
whteWvIudKTGID1szZ/RcItDnG+vrVlAG5FsZ9EXYByxrypiJoLUU3jF3iJm
G8+mi2Ef5TiPEe1kY99VR5jcfxJMUweywTHX4RocrmhxvXtAbkpxKjM8hqdf
1e70B64apbl6ZFTP9uinS+yL9BvXdDPp9EYORzzqfHSOKaZS+TbvXs06E9ND
oDabv7mZRT2EC4R7dIRLTlrfMxwYrWavOP8W8BUr+3waXjo0E5fWsV6S+td7
frPvkuiBiPGeOeWSrQvrPO/Al/ZiFwC128b/0Z0mcb5FR5OpDwOJX8OkoZsV
kLchVhLdzI9Eo9JF8vTK+Ok756c5GtYhk3A5QSxnRyQJVs9oZQQ9sMjcr+9S
XU14Q7o9rkwUtJF7Ig0EsgdHpjadV+/hL3D11cSakdQMPO5BS53l+vmooxc3
lAmuHad/gN8elhQE2YpvGLOqM9Y4EEpUcIKKWMSVyVc4cXP8+xI+npGyX+CK
GQewwcvDYjKQyzJe8n/8LNvb+2QxF8lg70CpT/Ru5N82SfDJBVvM27yaCXDx
C/1OI0/94FI/u9/1f4/QkulgZIchcY0t4uehCqGdXz33BEwUZPKkGb06gwyM
VyboB07Zj1xpC9UZGUKxrYndWHAtku4ztQX7gbQZM4LWGLdZhA7M3014DjKC
/x4J0sB6OSsTa2GGcAWZ6mmsBmOmKwyYs2+WWHlQ/4MEA0aB/+ARxtQjNYx+
suvj34BARXCUwocQTKh9aDBVHvzz2zSVBnFWj4l2nmTSkocqmZYhqSB3ZrTH
g00HMMzO2uX5d32zsXz8Rn825xTTmN9ixj122wNZT+NbNrTZpI37dPhtf9K7
wBNbX5bQ49ru9rk0hcV/SWRmWjt0ktW9aZ3hpkM+rcoln097M3kgpMb2bo3C
XMKLi5unYZl9mnJbEWnzHWbOIcIqteanAHuj391fTqFOgOXNONQFAYwfZJgY
Q5j1TBAX6BRoyqpzeaNNXm6t4SvxCXCYR4/XYb5xKVZTI1lUB1j65e/CsonR
NAzbF9Xkon6R0G4mxl9iLNKYRI0TbR7oRxW5zgBvs2kqzkCtxFAntUaENmWd
ka+EG5PAM8paD9gdqIROrHLgHuWkqIJhdlCjqgRw39V+0CGA9FJ2xsSDf/rn
ccDUk1CzUPCAbesigc5jXXMqPVDHKdBaGFDzMt0v1kWsn+Qwz8bIsVMsxfCr
IHWrNAZ/Rkz//qA4XGx3/ICE3PwDWBRtKecj1c8dTn2Je1XJjk+jZhtkDfXz
U+vn8DMkWXlKsUn7VslRYPImkG/wj38fKAgtmvupYxm0TooTqFhfrMtjD7s1
t4X8V1pDSj5O2Vtl/7sqbgAtUIKWJlds7eOZGySUsKFzB9LMl7ym2fwezMvO
u7BTqFiL2mDAQ8do3BWOsZNxlFBEawqoARGrVqkV3CZxOF9UfaFaQDI1qeHe
tnTbkxGzoT6Dj7xxP417ggQRARUrQMWBgf7WivVKXygZz6ssvNPSB1TvzWGO
HMT8P9CzQai3LUOfzm3ALASSGe9AqJswEAqh4SLb+uo0thoyWCRzvp7pYkcH
hO52wB65Pg0PLk6IgpMeOplFtEZcyh7mdTYOZB5ouq9xQVVKJRC6s5Vo8gmE
Fg1BChxj5GNpoNuLLKqkmJE9srwBZ9kbwJTQVrMGXlOxNRiAgXfc51w507B2
yDY1Wap3L7MTxfd9pfTJmj0HXRvTBg5+cShRfQP+mJjsod6NegexIdTziD/M
wQT5NgxFaAKW8HSSPYiLwNodN8NutybYXt27+rg7DAxbOS98yozv97PQH90C
nQn3pegou1ouB6lN2oQsDymeo4ZX+YCXrZWs3Rh6xWP9DB/IgpntL0wkFdZP
NAxwJsnflekcCylO5WuhjvXz4cZg6ohsenZ0cPAtzPzft3/JHHUqW47wbKhx
/mmLqh1Bk2SV6y0+yELBkgOEb2iovHmAwoEFaMlHZ3IG8yt3fe+L0tlCJuHd
kFO28MgRhAA+26+Bk6a4LIjjD7Ur0w9OPTm2Is8UQS8XI4dIpEHw0pXxTrIu
Fv+VW1xLssPg/K4wwfZFsSEJbQiY4uXvDXdXJXNN+aKPokx4mqlvsVJjYdFp
rTa/12GHq59XqjhcGI1sJW00gS1sSwWiU6er9LRLgA0PBduFuB7IW1tE8VYK
Jthz85YNtFv3jLv/cSIr7L0w9HFC5KKiQD118ZPWjRa/bNJqs2CHBIM3/NLs
F27tX4aS61oyC/H/VOx9K1B+9xs9ygnyNZXpguHCFbdeFaVqq6RuQyU6CTiP
zia9AJMcz/Xvwddf/cqyBGHVXOgYUpabyYgIMvYrhzGBtuvHpFKa0BFBcYZO
6nO6ruhZ9qMFoASWmx3KeZ6S8PyWqYxzvxQpuEVFNVwOeX4u9z6DpgAOKWJD
AJQf7gwUFL+Qo++qaWIBLxYe2UJzVfE1bmkoYS29yQ5RWc4YHfm4w4ur2ib9
uPVWTG0WHf7qZI1TEAyCjfMOz4tHGhwcEoFoGT8XCrhpZxttLCUKyiLnf7DS
WIYjNxcqbNO0Wy93LnXgYgJEzgQQTPznznR4qzLaI9ItWgg0RjzDFKPXkU52
EbzwbV+0eBdc97jqr+GKbD/KUvRaqxSkCjuruYME9ECatjc2Xn/DR63MXcm9
lbRh3wtauJS7nn9psqt4JdAuV+sBuhzAKAnOXe66Wqr0e+AtjocOoO1T4+iN
XRuAOoHKeKqhBkaCn22B98IavYlXSXuAayGGqep3kHJuNCFHrq7fwNgTQ0Fq
xGzWl8JaTXzm38bW0QBMhpa3iIOzoS/NOmjjxgTiXM3ZyUxYT5ShpLNdiOfw
YWJMPtiwoAuYOObaDPQlf6DmolhNY8az+XBtw6Pq8WHY4ike5aapvYghx+LQ
oehAOGGGF/aDYHgKc6n9HOMyadWb5ibL1n+F+4ut1DQDEH0l72vHLs4Q9hEs
dr3vVzLr9s/C3HvQfjB7FkqcnnIHlrN9r5Id6A8AMk+a+K2zH8VdTmd2QOC3
VAWnY3GVQdoJJTAiWWKHBDi8/J5+/mFcf43fBGBJT1WHbc83PcUBLQ//Ed14
6sh4icm6BAYE9FbG0bDhnYjcqKPNhJnC3g5sBP2J5L68jAS8DzAqR5S3wCeu
UzntmjjeeILqDmdrjPluICAI+Pf5q6Rh/a5ueu5x+18QbcPanNRPgYRFZaeQ
m/gDJi22xTwQe7v+pyG/d8+N6Z51wUNFUXhZB6b3E7TKfPPorM+ATfIce4cq
dvUsk40zbRqzztV0i5A52uigv2HFZIVBWLYYiIkcynWrgFddC3deQSNAXaJ9
eoG5daiCTxH11DwEWsttYOAnjpJ+hpUwAFXF+FqouHkaogtfTutOARGOcACQ
29mfxPB9ZZB7/fHLfCa0NFisO5IIlV0iu66NhGLoMqIUAe5Lo7GsXGzWBUEH
4uiCm1AUmrRbOS8pSr76de/a0EXXzFmHr7OYO9Gm7wYvZVN+JsLguyMTGdAM
m5Ip5xpsNQkqMZaOnRUZwbO/N0NA8/R7Jt+XRWzMgpOoHKjBYmm/6B/0/1Dy
xULA6uHvLdGqkDx9mM41I67DgCMLduIudyhLqL1jC9bdcIQHePUpfsO8222T
iOCwmHCFGhUiEflGGAL7QfZmSH4p8rTNFRvWp2nl6z6UYesUuH2I+bUQGmXj
WmJmMGHm2/DbIdbpMIdau4R1EgaF8nCmffhHOJz48x9zhWprQJWwp9maZsGh
jqFiGKDkS+CdwV/Qvo1S3Zv+sW5j3EiRuq32MrmX9VzCVYjScBkC+0tiNjy4
5lbxlTLBadvwBK0TLYh1b3i8IhjO5rZLtKh+0n/iyXeve6aiVLKuzrMPD78n
Ernl95K5y+CveE8YX3HZx0a3oKJtB0ycKebZIZerzWHO2eGNnbyha3SsymG9
3InLiWOd8853do1kXUtCwHlFcv95ds7gQ7/wQ2e9uwtDcCKRxUn40N/+u9QI
xO+Eko1bMjMV1cWa7jVJURy+59ICuppYAURC7O4j593ORB0DOxKFueuO4eX/
TvVS13bLJtbOsBNuvmcTyseJVhj6QD4yQ57/Umxd3nChtdbZgxJ4tmKQIqTi
eHqW32JXfCRW689OKMWcvkVzE7MI1aMADWsC/gKuVJ/BpLfkn8fZVbUEbGoo
Wt+uEbN9pcWKTr4bNNeqjZY2j++4vPGmSGBj6UYcati0HEk7ukrXcp3UAGYs
grObE8Ta0e5SccwfRTCfccW66C+tI9/YNuMKVo/tr60h+wMjTJkHRNYyJKvl
ZHwZShm+2R6EGCKn36pJ69/nRyLbaZegEf9GL6NMP93iC2DSN5nZKszl0BbN
tJmjG1eHIy4SW6ffxe3Y7SvsNZkgiKD/wbLLeYecO0BOHk/RH5nSmO77jCoQ
HSx6b4nZN1E1eDXgZh0FAFN6udG6lPffvQOPBQvcWGdsZcc4o/0/WwcqfLY5
pAG10Hv+Zkxt5VULHmwjLHp613tRywgqwJmdcQgv4/1y2HeM4BhzpGuvCxMO
ghgwCMM1qkKViUla1va3yZ+RtKqQKTIAxEw0hm0c7gQDl/WBPkPfCnLIStno
TP6kbiTi5QjukZxc2fyM3DAruxqmwfdyl8F9p/6QRZAkIrFrUoSWLjTR8Xr5
xEqbD4aWPj2XUIaBAzurSatwpB9chxwdSNSWJ0C/DsOPoPrT3Z+aqvjMo/8L
QdnTh7RjhhTizs/DS5pfkMkOPCV6UPXRFYGJON3i0WOPW91pDTMGuoJMm8Yz
EtiJ0ec1fIVJjnDOhx+DugYcw5FtlZsIs8RK66yYVcfmTZjXHyEZIgA/CYYZ
CzUBcBI8t2C+CRk/7PsmznFCngdjQYkfFtu/yFdtLYPokY9v0vMgWtCOX4w4
RBOCjpVqH3ly0N/p6Atmhl7sMn4vh7y/IVIV81ughnoyuLeg2vklidr73Ipp
naWEwcVbj14W1Zq2mV57N2fDUeAiZodHUwQGX/syY/lKakBApIIe0Kl6lSsu
1HEZRllSnHcAsFEJ8YMEyuGapDUMw7x+7Bs0kz+JyV21LcthyQ5R3bcKr1d1
erGuJjJnyCp0jUzzjNzcaDx6yGoaDEe2PwlkTDvUZfKoT+HWl8zVurJDgXyH
SrJsDRS6efnRRAEF+CSrm6sHQN3eQiXK89QEXAjQHMpaQQx1PxcwbAlBRpUf
krNi6wrL6XNrAke6g4vM/hPz0VHYCKOgp9d+6zWaIpOeUxHM5maZTlUSu9/p
d1aIGKWj+jK4e+50AmcfoYDBD45PTrVpu+8yoJa8MGPIdiaeu82fVduQ3NXZ
FsSDKrBtvvCOAelzNPa6pdxqjp8cxDxhvO5lWM5NuFnFgMSaQQHYZKVFkzBs
4cm+Dghrbk9kKhRR8g0mxi4pyZeRW89f0CRay2X3oS/eTo2Hw0oNUrZtxDrW
Wc+A8ouIxIaQxipcbnjiMbq/86j/jBVgOwiTMqMlkUjRK8EhrfRDYa86CP+H
YegOpx2c7ufvkkHGk8J5JnuZKGAhCZBIMx0aEO3RU3Jmep8l5Mq7pp0xfDr6
K4oMshnly9vHhnYGkx65QZxl8mV+DNGP61agKqxSp4nhvZ8SFTvDf0WOTCkO
JVEjuN/LIBpDG5uqaWoSKtLGE2dGUiRw8+yq3vkcpY5wDNYdrxfl3GwqbBmX
Kh8ZG8+98YThJWJOT55/s6DSmYmGl4oMJPl57pIKu+8YGyTKJvna25m4XBYI
Yh3PthO1yswTcmwX4dOxEUFUQFBrwXgMSV4cUaxkJmzM7l2Q8KMOBCbFSqMj
cHg7Czl0CwXc/8atl6+PacCcLFWsu2g1+nnFHAPFoFkhf/mWq+z1jE6SR8vN
4yMdQWIOy+tCRasdraU+7eDiTwi8GMIocFafu/9ASh36b0MR25u4cydHumaw
nka5RYrtivTvLt+35OwMVmg5mH60S7T6jPvJ/Om2QQnIIUDO6iqSq4yM3z0u
3I1mhcB4tDWIOxerKcSF6rHb4Oe1b5EomuEGNFcJ4qXvJc9IYUmoIxsI5Low
2Q3GXCpOELppuHol2bmZ59ixS8DbKs47MjlcQ1J2CAe+YQ4zqrc9/gUiRYoW
P2/o2592YX6vqFI3usEmrshVKbMwfLC41lLQmxZL1ua8H0JPrIb54onkWz9G
0ubLqZSGUvacTeB64i+sjjJkyLKfmgaHIq5rF12+X//XTeeLVmIgX3ScvOsV
ZND/NxfEnnDybyzs5h8YSIk70x2XcpqQkFzJPq2gKF8Wz8/F4tEKGbdN59p2
YPaXmUz7oQDQ0F4dRrOkCz3ddSR53Lrj8/C6F/YygZSvOvrnje8+q1jJryUO
Gzs7hsNRfRzh0DnqUEZk0J0PECU8Psy3AMumhABxphCNLkFF29bmT4mrmpaL
/leqw3yBsxRDYVJb9/gkp5Klk6xURqK35p7NoKXMEaHQPNracHIvKymj78Hn
QFs5EhvSrtNiKuLn1YUqe4PbodNxwdJD+J1xmu4k9+T5KofdTmMm+S6pIxSk
i+l7mPGGNjSF86b3atCmDcLtPVagVyW2wlVX4101FwkdLG3e4s4NRzIvJAif
tazaLUMZHCdJZAHb7rmFvEOa/8/Cvg9W2B5F7x9U+TF1ImAMcgi1PzuFkPu0
8Q/Mk176or1Yp0+ub/z1c7+C2wq1nMRCZKrpltQnblQA7uAxjOfwqhdywSB2
09+5Zok+gPtYqUlFZlgRsmEoYg+vLsvsexR7guq84oVDeT0J5G28/fd8n5eM
a6V61QeHvJ2h4/3yL3/0si5dpYXpNJ5NTIL9cWedBKGzh4ZRUTt+BkkYlOHt
dxpJ4MOL9YSRT/atpRb7qLQ3ZJGMxlvyVBrh1QcOtfYRn+pJDnziwSOLiPtb
p3V08aXWtrnMzaeDB1nOiLU3zFWG9RdZvZ1zMchWNqulKyDZnFEvIiJzvOUu
EVfiFX3u6d0qviT/0EHiXMm9eSkWpIZ1arr84B5SCHcd/RGZQ7qQI9K/16s3
O1t5u37Z4vqdxv9yK8KsKt+vM75OJ7FjErtNp3Rh41g7u+cHzWBECmHhtH0f
UmclQeI4gmzJyhTLnZRRdofFoNcBDJ1pVEpk0sEspjW83MVHYHRepCPZ41H2
mobT69EgI5JNxMRXqPX5Pi1l9XYXdXgkiZGlQoSmUpyyykLhT1CgiauhWgGR
KWp+N6R7Vj//0cVKn4gsoXq/fPoiVj1LBuPBo9nyi3dlSfwVDclGdoWXQBOO
3Z8KTlthmZDsNxDVgFsoDhxJqaxQw7gJeVjV2ajwME7udduGx/ZDfg0mvAz8
BrC++UhQR0JnBBWGgY3htft9kjCr7lgK546K8TNA91RsilIiZ3qQT56H0Kdo
uRbhUkQkaFiPzq5fjyUx6FJwIbM852g8SJN5jmej/xU8pmCvWoqT3UH+3U6k
PDUWh77HbaSOalA8v87bgCDRAvfkGIzDwYVlZoV7S5tcBL3weOjIbJEdVho1
HXX8/+b0kWILeT1wWRl3szgbY/RaScSuWKj/azKaAOjCZNh2JQf1v4XfLIGy
C7d+3eCKhtaUxXwtmYBcOzNAziXWkR6RAYtIYMBi3gfaiqZ0H/o8f/1hFTr3
9+eovkdHRyHa6RgXFI308u5a464AcVMQ1VyKPB5gIrn9b0X0d8V4TkXXiyZQ
WPrpoQq7cbQ4frCVAHDXKmaAdSdK20wF6RhGWDbyOI8JkL8lXTHD3DiXZ16k
gvxKkez2OXzFMgGwd8UDunCz6MFFrGboaRazHsf96qI6mOjWbhxkCnp61f0b
OnPObiPg9mpkTpmzumWcAyEju0jZqWZ1+Orxt0CFlzmvvtOfG8TYJi6Gv16r
T06Ezr3SdbMIDrwnyQVArdFbDlCSypjdvtNyER1plxfvBgeBkhOPoKVWavjW
MRIuT0VsSe2Qc3ffL7IPZnVl5eLmketyM1AmHRcwVDi/gIreVlcTsH1hCykm
EPDu3rJu1eNNSgL3JbHtWeNmZJZyh2NQCAx7F8ZKOtGKlxqQFU7wR+LW6qko
8Bn/V/fNHQfi1o8DYfKruSe6yqbaTMTf5NFvjBb1l3+H5OAThUW9XujcXtF5
LoLAqkW9wzBIcDhmLwF7/9wpuK6MyOnJ86ADZZeKzqSqI0E04LkLuAxQkg5F
T2eRAtmzV3waoHZ+FbCPWaVxwQIY7O19srJfQmOy1+idIZJ/HrZoveIhDt/1
Ej1Rel1yu/enzEobaNkab3yE+D/RN6nagJiJAy3S2u2Dnx6S+9YmCHXAqEJb
+dhc9cfehzY91BCTD5Nv0eGAIYh14V2kSPdlEWqZsagjjI0COl33Fry7zboz
qmpPzHBh4FLIykQjCXHdgPdUU+sDvwDVnyo7vNiWmac2kL+0gWfWyAtoGoQi
P1B3Cet93tvwqMqYLQrQPL2JGjqtmVm14aPSncqjG0Bew+ib2Of8bxQzNhhr
73DGogIntxil4jywnZjfWBejdAuCg0urM/G5561F4XEV2DQyfdNjGO5jvG6+
NwsO132BGQDq3zrKv5OeSq324hTpOClPvPG9IRSFoQhPyG1VPjGhUPk8oN65
cnOJT4YPgJPjtqytnE29E3Tsy5jwijkk7LXeClb5+Gw8RSIOQS1QN4L6/8Ab
yIN45b8qeVM4Cd8Xi5wtdbXUBDwQOEOy/yVdObO5Wg7sVpHoGJzYUHlChwMX
ow/ruwK/1QQU7iT+QkAh1wdXCXJI/FoZTNnax1cbus5Yp4/pRalVmLsU0Isa
T0EEPUT1si6oaL3DB6ue+me9T0DMAi3t+rkAzA1tj0lY02SNg+j3eWRMLJt/
NPXqE7EYRB/5QF4o2iWKE/+1xVvsx8ati3NCdIyArj6GkaPTUzgp7Zrbep+u
IC+Su5eS1FktUoU9xUpRgR53W768eKhDmD74SXvsMQ1i9zePY0VTeXzlgm2L
daNjQ7S8Pc7SkUO1NpldrWA3NAp3rw4zH3MBXQQ2eMA60f+mgEWLF/Z+HBPk
j0WjCvzk/kULC0IGb7TLHsb2QAV6XzPqGIlzugJe3QqNwKniyKqfuwNWj2f3
8fX4bjsyu4fQcEkWDpnGy/jhnMroZNrorAqZw3nEQpqITpk4irOaylaF7jut
idjRncUcm8+Yvsa4BEm6wnS/JpzWBD/3w7MCGXKxaq2RXjXXD6g4XnxegVrJ
Jvb6Lq3SAhJ9DrPP9+NU+PcAxe930P3wXmpArcrZgFD+f3IzAZhmgPmwvMrJ
L5Uj9zrV7ztwDQ2pjaY6JeErhVBvHDEDN1hPO3/jRv3anne3yVhRwx6MnOr9
/ukezNBcr0fKaNoUZLNurNjYA+uS7YmQpMyCutdtt8Rey1hFSXhsL9Pso4om
M1ip+LXXYcFOX6D/EWYHKdFWKhInZluV7MCHYDn8gKxGmlU2sAoketnfk1Wb
cy+Xf5YkmvxWybQbstc9RkXcPv1t9eO/IgHZw/Bf2IMuP8zAxqOBa8IyQcxr
IPtZ7qW1Nu4zsVQr5FBDghbIgB65btInMJEqeVVoWuL8KC5qqwIpZRWPFdMj
eULrPKIVqfIXPSZsmMbe7GlqoziTmkK0FqJ1tRdpOJMHYnnUWUaw9/VAVNVl
NkbFAW1I3elj+H98sO9il4NWH2trgHLD/1FY98dhSmuumaWMdIA3KJpCu/hB
Plc03lk8gxed4HQ6dOqkijp23wACsZRDGjn5Y//Fsy5Pjx9xbttHaR0684S+
Ug5nI+vQvG3nKzj9TTq05iiZQ5uwBzcokNbF4tKYnrRU5wNsdk2Yn7u7mHoA
wYjcdA3r+GTvK8dT1NtqopFGWqpHux9bjT6D8bv9z4A29VRGrv6eb74J2DKS
Nl9X2Qv8VSECnVkL/zhNgZjdGXlyWIV8cyehIYKuU6r5OVS8xNOL/ykmBA4l
64R2obtNYhun8B0H+wJz0BsGKDSFIozoBtlkhqkiGxu2OxMYve5vFAs/Z8N/
sDNeS07DX9UHcy3AeRTThX7NkUZwvZFWiQWupxse9keTQG+gqltjOlAznNjt
juXB7+lyGjdGy0SdlNAqCvDGmadmhIcZ7ZHtJJJn3U2zfmyjTKu/H4vseZR9
1YDTLbqhuugQ5rEFGQ2yJru7LsdiEXA1i1LJRc3XMyCmsNG20MmZirMDzz+t
CAFSqRnxb/tmYQ2PL97MuHrqIhSXs3K1X/6oc351QTtxVCDgosbP9uPzR2PM
DF2PyqZlZ78FM/FMVlCU0smVbubz73lyvoyliGBOsRAZCmR8lMb7RYDqXn3f
8uXn5P5k8+9c37GbhPSylVXbDpudGPenZhoe+LRCS16M9netUDkGqrNDUzVt
fQHDxSSllfmjApesoDsk8HPJcUU6W94eiXuJUNrZxihTj74hV0yJvljiEXPo
xEiWLoUXJc+TWhwKtYfEx9FcInstIA25II8vSXN6eyQomb4PniMO/1sdkC9h
neFBqqvBBoo7kMo4taKS5We9VhGgdFKjjdfrG2STnNxAXvdJapi4/UPKULRA
ZiRbk+RVM7jddJtWbvBxJdUbiH1RKzChSujxHGd40cS92ANGDbM0UUEBThd1
dAQM+qCliUAsEltbzr85amucC4d1cw258m2FWTDuSFjBGcTf61WCq6x7joBJ
3IwE3m1+Bn6Mv6j520SQQrDDdE48JCmriBfVf3DS8G2fUB85pX0LFvv81e+p
OGqVE1cq10jAt/6+6wDItRGXAbqNUDVRBD1YbgrcWSdpiFogk3j+0tnFZpZa
bpwktBN8Q72ofc88Za00HnndgN2OPnF0E8st83Zw1spyTiysyEAuGuXBbkul
tO43zTp49UUWNuHJ3F05h7uB5XD1ekrxKkrvnhf6VoUqISvCTnwuhEJqBQ3a
mVQVK0rTn56hWnplptJQ728t6X38y/gPIbFZKNyYQiBUXri3jMlbV/CNjaTH
iFE6E5B8C8cZmHGs/TvqWf6b/OK1Ri0u0HglmkqpJt6ToHDdwAfXISL5yVHS
MJtKtFOzU/t+R70PiOUCsYWW2DXl0ymbx0lab5YhIWCifiv3tpH5HdP3XxyJ
L8WKRtN2+a5xjL6/9Mh4Sl3Yq/5UoYKrZx7fF/2GPQJVenr95PcJ9QOwM2ZN
/3XelS5jERYVdjkKYQgiAkUHoUNihi+OoqkfXrZkEnLjIMKyYxulscYvFJSv
emWyiAuqMakWb1nyaxDlTaIV/XRwQr9XoV2lQr2fCttRJe8TUYLz69BzZ1/t
Ze0hpLzZLV9tAPnCz3nIj13+kehNdS7UdZJ4soGCbXLzfQhHe16+1Bm0KQeU
gT34/IsZ54wWiWgAFVyCThWjrDA99SkP1YGxNBqXvFbWlkZJ/ivV5/PZ7NKq
DwfTf1DG8jlnsx8xPO5GXhXjvZU/fNbUsmPYxSWMo07W+XqKKJow30PmydSZ
dnFX0JQCq2MJNAPg21bowkVFgyqxD1dukxcSsWFlzoZu2lpw87uadrD75Us+
RgbEhaChbHhPJ6aMYgGRWRnvLOVwPXwP0ZKxhEmFk82jL8Dtz9yp96SICVZa
HeDBKxnXovZccbkvPbo2odWGs78cJ+YAKjg8Bj+NZpQ9R8DxPLK5jbDgik2Z
BmqD4fQzJffNkhIIOYooNTtTShXK5mXFOGjtlB0ZRVRGbQzD3EkBJeGcwXJr
DXs24sATn8O35/UO+ak+M5/PZgCHBl3/IlPrFFgLUKMZ0bZko6f7OFvAHSRD
fzGGJcgAzeNVGq61ugHUY1euGDqUcIDF39bB52W5ZLtyR9Js7G4v/2JTC8mE
p6g29SFSBaWgWlSjKVXoABqn/Gap4B2zR4nEgQK7++pUxBxOI5nabvDL1vno
60VIEtoWncdzVJ3OwD6EoOqXVSzHYWCd1/sQsuOFb0UgacFPiORg+3MWLEfF
wVhceaprTK7+BxMb4YWAB5SCQS4n3sdIU5SX0J4gRWnmhIq8jtFvWijb+xmb
ysxxU0KOKS8QPKgRRfFi4ieDh0N6NdxGj1XNJaNGHEbyFZDpU4h+l5KiO6bk
3TlveIeNKsilyfvYtu6ZaySsYnxA5KgfGzKaQXS62DAPVzd1JFOzt7Zw5QEC
4UaorDLygCPKQobpc0VesSzjkN4tpdwnm5IfkbAb/rpNB1CpeyxN9lWg4KPi
d4vh6khzd3fMhnqfPPzzB7OKQ1f/yEtGmHCvXXrJeF2Ed7DzfONA4Vm0fMTT
Z8uxzG4j/zrO14ZyruT0/mWxLoGNpkmQERZnn3pfz49k7rajp3nsnV5Y8/lc
lNgskQJYr9rRG6E0DVmIoO3nOrYdncZUg/y6clQDJqM/bMfzaH2ENT4aDqE9
zeUhlLRV9cdjv4dfw3Vjqm/D6NwOrwBuFTqKFMt6AoLy11Ibq4a3zYz4FuNl
NG1J5EL0zQTpL2uSOjWkgWRDWAB/0I9nZViTavo5isByb8DfSjXfaclIbRvz
3VQdK+5BOQ67v2EMthfAxFa8B2h4aa76cdivXKnf9QzjlHL+mtx9oyYqNLgU
TjcnMMpbIx27Tq+7ExWlrwn1rbyVxwo41KGR5LEQe2ZehrQqZPQOwpEOhGUY
VzeQzRpx1n8AruvkX+R0j+DoRdbVHNvApPn3mFtxrXl93efiJHfZAoOTMhFB
y6WW/cCQda0sSqnINB6/n4x16mfuBhIp81sodG+CM8O04lftlC28l5idObWy
vfuasoVTITjWFGklBqj8EIFmoLoWye6uXcx01CWgSVpoCKD064SKd90XQsPr
t0Q+8H3wqJsh3GW8D/Qtoult/UWCJIvFMCMQsRgyDtrEe+Sw6ya8Lp3iCw2p
zB4hXejEvhJLicGJkxq3NjsUMlBgCB5VTXd1nEhQk8tcgg1MowTMC+zcqa+a
NHoZf1MQqVO5Q/rl+PrFIPEWJAtrOHMBLtKlFxnf9ArWlist97Bk0PpD2/zw
46BBPVs0wtfSWQnmMt9AgvtJC8p9HKgjR4mptH6qHphbRodgLHPgozl9Tku/
uuTBvm5wtnPEicVl3RhFXs6fRK5aficjxg9EGg9hhC7UijQlhJ0jfvYLJq+c
9RQ9eQi0FEk+oJ8HuMMdJbRz1j2x7oLkFvwC+kausAc/6/qNshjuaTi7oTH+
QgvZOFsnpmLMaD4nF6OXsWtdKVpM2gXZ95kq2563Wr7AbzJ1TiWB6d2gEkTR
NpLxheu/Ji93GD+bQL0rq7zEPdIglVncdOGfp8DKyWr5E1duOKp4g9ArZ2tW
zlxIl9Z/+Ycvne/IyjX3e+DKD5dz1ZaEut/CzFAS3TsLYjG30QYH6Nuar3KM
eLPSoYs6SMGXxbIU6Ef/P24pfbCvQa7t5Lect/q+27hlbhS30VtT4j2YVWup
SHIHops2UwwlmSHnWAuzyGYHw4aAU2Iz6L4oBGCw8vFC6x69gJQaBPsYrcn7
iw8HNY0tAc2FhaONAuqvdwErrLMAYQjKNMtKMofouQdNSmYu2RcxR03IqINU
7u5wpelOBfinogrhQRgEVjvkhYirTPZEVpFpLTsMU6it2+7nw9ghkmTjA+Ei
wCBvAOEom3BagCyMi9qnjpKhaeNp3N9tJ2DQOLN1595OD8GTnnawB6lAZ5HF
U3RQ2nbCPnMHqMP/ZW8+u8J/5Hj2H4s7lFOppY8dx5DBC38puFgrdjRPyGAK
cJbdo9FVK7k+qbIveKHVPKjZJdtRKJunYquV2o6rhVMhylA9wQptbu01BycE
uN+eV33AyFvB1OX0W2P6AoWSSA9d85ckEDCJCnlnn8y2wp7s/eYCiEkqtTLL
f4nHw/ZM9VxB7zcHmM9gkpL5RaF6h/Zc68Q6jfmKlvsI63IJBcoxtM9h+lUM
/62pTEDYoaqaXWQiPuqV/9YkeBiCOoVdEA2tyNE7EjpbWBPizY9PZk4gKlxH
DquermMeBhfC/4rjTkU/ORL2RUdB2ABePG37uNiWXSOGItnKURgV4OJZGq2O
1BF/0q8bNwaF5IGOjUIUOU/Q8bKnKIcGAFtytYKOT4kcbAYfJXu3ExDBn61d
Xu3KwvyGLmCcVVWUMnolytCINZKA0Yjov9/25hAwr/ef2Hf07fv2aOlPknSL
Lx9R6fkz9wTPuV3/gwWy/mXSitzZWOCFDJhVJx9D6FFnpkZ305RjGQTmbE5c
3xkORqDQlDiiUTMrztoHh3p9qn931XQkjp23m8qNyJryyQQE1tzJ/gyCaErM
4nrNp1kbTNA9vFk5vpJQrh42HMXieN1V4A7nFWCG+RKpOcDrQpbbY6jxh2jo
LqD+OF/EtIGR6+v06gEmj+yeXAv1qsa9T1dvHKlG9XeFWtTHoXYmJfmvqet1
/Q5jfaReB8wFAuzcZc3r7r46rG4hq+DMcc0RK36P9fxbBrLHc8TTFQyMdIyV
O2csMnjafd/WUL6Z6fPqwa1CZnNi680igU8rso6U0gP/bq8n+7HEjaqsHh52
0LLHFgNfw+YxMaffegc9m9Okv8HVK6hXDUuuBdw2iCaBGig5P9Mujd3wUfuk
rEh/KcXYlBkQRDrw5qATjnXiXpVcLc8iAFkdkmjLyNa/9bKTVc8uucmrkxa3
M6g9fGa0ndCW1QlzWg+4VrSasdTNk8z2QpemBQlBhTgdf61B4npRGu0W+ZGB
evLrbP35X6TIcJOmn9AUGLnledtvVIJ9LTNqP7b/2/jKMSyIBA2BD0RDbgSt
2a2oN5pCXRmzWz1NfQzpbj46TLWvoSlvnQ97EHadTTDO7aGE/dYOpzmbGhT1
dqshPlPbT6eiC2j1TFd4RH72iBWDB/lvy4yiZEIlizQbPBYOAmFwRrrNJI/b
iQb7/vUjYAKE0IbDP9d3Vz7989xUzHrpupjkUH8/+3ZhE6NH5sM5WOoGadhv
FDblh/HrcSZLFSv3LDiEpHi/0QQdJcfNl+zBvkGf/mTysMuroO9zAEO3BlFo
qq63TG34gw0pghIJsatmFWtsdQoE41AV/H9niNb+kRLOM4JGpkX6Ji8U8vZI
iu/TkgXSrLHo1izkA1ugJejRE+Q1wgVN386zWNraKlXQJkK2WK5EaLh0vhdY
J9yxCvDWMIgEZLAVkjoquqLHi1DJFPVs2c3xTWaC6+ZeLkGYz2zZo2yfViA2
IK2uIWOOoESI9Oyld0pcWDIabvw/ivggoGmugrVTY2w62OVUDLPbUC8gIU7u
SmQnZohUBOi+WG2AJHGezme9YqVWm4BAR/o16qfmwt386iMjM2C8qxMjWqIv
ZAUeB+88Iz4+qn2nz4D5FxQbnIHuru7n90fdMDvOnX0cVRL/9s+PojB3ffRS
EYTuPwplOJZ2PKHHvpU1jtzyAYu3r0cEyxkC2BedDUsy19VJm2mf059ZlUPB
c2FNPEGsJNI0zULZ/GMLOp+oLl+5kDv3Dtw1JBcWOVEdMhJK/flWvoEItAxm
GdoL+I3A/XCFcRfoZOET5NR/ZzDP/wyeLgF8OOEvXKc448zsukL1CnFKd5DS
ApEwljgu6DNUpaGy9KSS8ZURoESX1nRuW8qZcQf4DKAZAZnICSQVq6nXtVb6
g2O3EhDeg4WDV8aPgSLDPx8w5o3bh1u2iJjD0ShbOlXBw3z2AkyZ0YG6NhH+
8Mqlm6VmeCyHlu2q5sQsHKWDtPAQeKAbpBfXa1w6pvw9qeE/6hUx4CC5f38z
GyzuQahKCcKKXh/BCZA8ABPBta2VkabI5iLwvqAsfKTLlKQCyVRdgK5a1o7b
aIVXtMWGe3sdTz6MKWhig+EI7yrE2eGwG7dEN4GnYMHH/GrVgm5t8NlJi8IF
ilY35x+mqvosxAiqqh/6ODzrG/NHPsCFLtIDzPVAzoUrjFpW8ui0TlCOZCSC
oj3YI7vUViOTYQGNTbXiK1aZJOur69cpAAt9v8RX2p4N0kk3knrFO4i7maa9
6YzPCvezK/GaLU8NXOsUfA+JRCF9jGa34x0eu5YPOXLJmgVfN82dLix2jzrb
3p57aJhYOJbT0D+69BrGRjlyFNBT9V+Im+gKyPMHTuX6SBLbY4rcT017pmog
/21/8i7EngtVZrHU2+o6655P2S3NnLFF65rhRxX1lwiK7vHRKbPGvh9KsBY2
+AmWEcELVsMyJjA4jP983xzLuoLtUJuGPXTomA/Tpk4J/jKldsucnFCVD6aY
m11VMh66akKEebnjDM41civShaTsLAymxDL+ai2iBomlyEe5R3U01AxZIr7G
imcA4IjFXN/vDNVR+CxRBrp6bU3MJvxJRInivhWG19BPbojs2VzZYqk7sxvS
M30em8zLVD2n+n773kcgOa3v/QQQslKb9s6NEMDmR20OWXDZitcUOT2zP3LT
qEUtegPt1FE9pd9nz6EzQMCQrqcaajf98YJPoiJRDe2T1uwR5H1SQAL30YPH
+I3wZ1wqQeUgGC7dOt8fHI6KVcbGyqsOwC4lNZCGopnPnKzdEmOfeDKhsJNE
NLOJCIR30RB1u+9r3BRXpvM5a4FE2/Ry7FHD2AenvRAZ8A2e2y9qwxWzmsTk
5yxp9VhoEfk12YxvFmULkl3yAa6JJZGreU2NBPHnC5WRXWKfQR1jJhzWYuLu
wpaOW1TED1kjNFZ9u4EFvc3IQNJMwBfF45/M35ZGm8yx8tL9D3ZxDKU81sJB
q7c8khAA1/YOqZHhWHPDUD5uTQYLUYETHU8qLRoK7ocnAfqKKGpNC39MmrDa
heztuewh+wPMCendpUVxOxrjTiWS8i3Ox/Qy8QaErb4p/HdhdJCUTKATcH3c
e7OIj8gLKcfzFcw9FbF55owX6CoAGQWo2yiiKli3yvp9G2H6NxZlFtKDzmxb
ihuc1bYiWPQkcHDIELgvf1ZTqapQ2uTadnsP3D0Qy2CnVKmJOrv8ug8cphS0
/ZGJuigeqvO+sqr5QMjz3H2m+jhtT3/T+YEaB0AtavKe7Hygk03Cgbh5iBHT
adBZyf3nTBg9xxuzKZP/09i7GsgFKX+HWfin/WNNSwdwJjOfaOE3LOyMfl+7
m5U6KOrzfomSiMjS1imTga2+O+4Z9KUdLF5ut3uN5J6Phq+afJndvDu+tXCX
dtW0uz2VqrAHtWVcOZzhAWysajeCixBIvgqwidtKvydyeCzcPFKYnPP035pc
nkI7urrDEH4qwCvVeL5uEp0aQ7QvGIUzALylLPnGnYtc96nszrst44PKeW0Y
79lBBnrEM7XauvyN8ijq/IrphnCU5kabsSfUAhseodgmqOPnZu3cgII2DXPZ
gTxuG48rMyR/TQYZ3aK2to1vZuJ484g+2WqXeQj1wJ1p3Y/fjEHoO9OFE54e
lnYo4rx4piXqUgTtxUlsafOIyR+xtDvVu5HyE3VR2C89kgD4YC3U6lltbvlM
QrOixHBSJQtR9sdhBOgjZxn5g6x3nK+hhkHMJXioV2HxinZXscxjiEchz5q5
i/+A6j6dur0137pqO0wk3fzq+mAIKiGCddwyEsdv8F3nEZZj7hpHC+CUOfb1
d/v1LuePRfV3pKuHqUBFEhS3eJOkSUY8XLcUCvMjkM8S1ZFG0/4uNccy7Jrc
iOnH1mBXE3nVj2PMwSMzz48yE+hZi2JNqRnVVMfi4zmix816WZTa4E/XrBxU
Oj0H8n/wU11aNgYK8q2bV2vOF5mZIo8j6F0XgQ/Xj+b8JvMytVz6JTmFgIrU
Mziv8qz/9p4ppa2Bful5ldP2XR47ICTwMmlAsxbOp54CeNa7K98F1kvInhcu
SU4ODjhE2Bter8qXfRfiHqRyw2v9RaUyg2sxWodc81jQN2Lfjvg58hSBfyUh
YdeEHv8RsowJ8f+xzspIMH6l74Wf7I1IuvMoo0Pig07RgVqPd8KK+/PEh567
BWqMQIH/WPo2Wfw4CM/Z3TI/aFs4U1G0R6O5gyDIvCAhLyTR6kZg1afEtPbV
Beee/EpiXJ+q5/acWx02uVVBMWdXEKDiCWpK+LJy6+C3+L3mUoiwdmDlr2OD
i/2BSqkmTPm6XCYJOuYRv6vis5nk+wxJ/8eng3BN+pctVkiErnk2yLkdmo2u
K1gygZn+oRh/7Ym3TMgnbOKgDB/i/PpyoSVbI2tAA9wxHkCisXY3okqaR8yf
hgIoYYd5IxngUifHBKiPEGz0lYlm0L+k0pbesgCnZKJ7/xK4a9JsiM8mXoWQ
zzcOGRfT9p9qD/N1x0M0JKPDN6BojmchmMrN0VEqsH1RWESgSkf19S1uxeKt
Ol9+cnFmkgWaMOUxid94rwLyQKX9noM4hByF58B/kU+JgW2mzzcE2wceKbAm
HQQV2O4eZLvgJNZ2VNvdGXH16ph90YYJKq5XBNKzLw6znrXqKBu4ovCV/dWS
3yjaA2X1EVk/KWNsbOuyU4lKTPyehdHs/iqb83uduDlHC+8Y8FZq8lT+z5kR
eEb6i/eHknxWDnuXJklQMsg8dzz2yVSnQSJrltQ60kO6N/rfUzLEd6Ge8Lrz
wJqVIYiCCAPwYK1fafDndx34gtERFvwKKGKdA1t77pWHuo+RQqpK+oH0hi+K
SDtJfEmKgcybBRcV/HiCRv5wyPKGHipK59Fsy2oMRsRhcATYFz6/7GT4PTOD
r/TPRnjdHm2gw8/gtR0PxBTsdkD8Fe0f50t61dWzZUYat7W5qRxBHPn0hJlo
ruQjBBWRVL3wiJpQS7tEBGXRUx0/+8bitrxR66uopaIufXCvCkXpOqdog/Aj
v5ApvzpxJ4Ye7qy4tJDFX0AMNF8S6vjbnYiQRquQV5v+zO7D8hyaCkTJ1ByH
rypsP4dz3s+WXBR3Fx758GT56hkVutvlOuDILpHcFNweap4OSbxwqeZwxTuF
NOfq1UVFZBdTZtJRsJEwPLurVkHvnVUXOpzWNjpIyeFbbAInd+1dYfAGwOl0
d40mRdgx2/ekwGb0Ms9TvRhk7lUk0wSb0jLwWtsDnzdJ+Oq5R2p1FwyGo/RX
AWNFTDCop1x9rJXtXvUPepBorQseOWpUVZNNrq8YJjBKIkespA2X/PNqfirp
GEVVlbAbOsJjA/4kQDUGIdlLTsFsUsaZKhfnqR1G/cFDgZW9t3O7zi5QMJCz
FPLNUphUhXkwTWMwxzFF2y6fQ4Kw/FWYguJkuahs2E3xWmG3rxfp/VvaN5PQ
GJThWrxqboCDpIoShFV+YwTPGa7p7zr/rJc0RZte8vnG5QqtDehMOwzSftJp
eJNnmac37/i4jQw+S1RQuXUEdMBXiCyXeprlu9rf9pUGPfQUrDttCF0lyR2g
WPlqSrfB+w5JqQqdTmZDQMN35JQDx8i6anRFlJsSsZjcCT4Asc1PLdgeQzhm
95upcjHAB+5vWX7z1qIsmPBXt9dmdWWuaHsw6TMTAWDOYWxo/cdZe6tWYdHA
77F66rTr5flBG4R24L/a+ijFUSA8tLXq/J8WP+oL90zJWccb3Swz9z2qehWv
tk6LuKXo4M6Kk/Ay5TcnrYYZ8Uo09g5xgi2oAK/shwhwUuu/CRz+nNjVjYvy
jH35OIELy1Kj4cU3CVHMSsGSy6Kh6dilcOjOnMZOhwsbwscut+Ro0AH8XHzj
T7/BDiZDdxVRtw+p5qWykDx4m6S74TwwFjk8bjKi8vSeQeh07IpZhdzKx+8v
NmmwDnS0EsTxPh1ezo30oihBG4vDdTpRvjCfhb3ssAcFnnK2IegdZIjvWC1m
5xadE28/YwWHGAerieljOWzela9WWPd8ZEEYohNBZ+lawyOxMuxHZciZpoAq
yasuPmEhEl+4sYrD0yX+19fc84o4QypCyJAU6NBXNWeWjeHG1vdWCE3NmiZ2
vAXNoPssGyIAFKqLQJ45JZKZYkJHC3MbCEwoVmZFkQOWSCJHne2Syd/fbnRd
p4p1SD5yFDpodDSPMEle+bFlYBo3Y3pLgjDwrDq2qhbxg2IbXKSR9f7LbdkG
NfX2N2JNk2By6HgCVYvrlk0XFc++IXhJAMnjUA3KRTwW5o+TVn2K7cUpgkah
3evosltuVNetopi/fC2guU25n8br80eB1lV4zSjaOKFMj81whDk9N8ZpHdR4
yMmsG6isEVzQttBiouiL8dPIh1lVxZPlvb8pY/LyXrEEsjdVquAwsgDkCEVs
TKawTz05n2IK7VmPBGhR7/8faKM3OfvOBP6kKCGzhNbXBtv2lqjj0uVyJMTV
1xSK7mE5cDhhf8Zqlb9nWc1g67XRRrns1ptRx6f+RTZriAyXhMAqJTL0qi1p
HXW1yi/DTVl2Ysn+bMknsZV/GVMIBT6fG2YReJswJFjilQgCg7tTexW0LJ9J
1nZpwWTSU1/ObJVW9EQDBtucH5cbOyzo+qUWer+Hq01Iw97XkyXGQeIgRZbJ
hnEftJYqjTRafS2X7X7LBbbDsaupqosbkeisM8kGH6AlbcH+LjzMC1sJ9PK9
9JRNCAmI43Jt5pI05Gay9nEI4aT0XqT2hzIg5AyuEq6D542BeKIMh1m8aYZZ
e6MRTh52d1RnsUb5EY89RuBGEGuTIYxkzMIAZwDzUeX4Msp4cBaFv1nUW5HS
groi+Kia/2FYv7jv659bOmLxX5cKtibL7M4CJsj7F8BEv9WzIAGnxOF0HwDv
n1nRUw656tYra7cQ+GCyPIOGnBfg0BJjeWe8KIDfXgjoducotiy6Qz6Qyf7P
7NfF505RQviunAX+1Ry6ymbAj9CGqAvAZy+dzeG8KjCNlcTFzcK/jiy6Q9Vi
dYqls+PdVRzvDJWcoCkMxSUOYoNBUYgeaYzI3Ay2BUysvOc0Xs3LnyJRVFWr
rxaSH5qFLtzbipFYvAoj0x5FXqYn4w+Y+jISFm1w01Z7vKrjktjmnk4z4S2W
tZAjwvf7720CtaM0SybrW9doGbeZWUZDc+hPekWKcXJwomUxc7e36qOr8AiM
ni1nkFbyx4SyeBtGS5Qi/zZDBSD+gY51+6PDTivJlKmNP8dzAtxKzgohAppX
9b0PXiABchmbZVN4NG3gyuRAcpevMuG/eddFcZpWZr0wqN1M3Y9rpMbKvq7v
69HL61TzwR8N4GplGUqSiCny3sUNfPuFfiWeK2mFhAMpwjjpV5kQLVQPNm2D
KikoIq0eikA0wHoG7xzvV8/GDDk8YoaFAMYRTOrG5mxZkWWKgmrfWq85JAhX
e4tAoYVRdhLvFxPNothT0gNVgvHl1QRrvIlIfwAso7WhPGzGjwwG2iVLrCD/
tx28T6HKQscURTT1eBXYSGiI9bKA51H3rLVGbPzZMgwD6z6/eDFeqQeZ2sgH
/jxOsX41Lc7iLdEzNNuY743xh5R4jmVWBfbKlk9DegmRh4C6/3w6TLHSS/S6
ApcgleAQ4u3Gw0KOwNETRtONyFIP3wx4jgLkPDfpR3wG3JAZsIIgZgyYAVYa
+UoRhp0CR7cCVBbneN01pi4Mrtyr22OYI4nGN7JCliamT3RLklvfUcmbSDv5
f+Vc5JULqHOaJgPZiKqKC0JUTF6eRfnEtfC08RTI80/8j2zOYWDRzw55xMRv
vSOq5fhemiQ41/x5KQfvpjJdM17BJSS8SHrkR/yrGZ0rd96Lw0Fs39NemjiB
PGx57ASFpDjJ2Jyd8y23PaneKUrgHotOoTeDggY15TwW6MgWmImZhJapdDlW
pIf9f5yTFnsi5FhmYoXMEPWTH8g46iQiEd8VqsY2Fma/wxeUuabgSK2MiSc8
8nqJMp1m4lGoI6RXLcNBFolU+y6tC7gevz5UAPaGP7zE8IHTFHRzLVavEQTN
a+r2ixg/j/52EKry51Wepv+8NCW90Uz2x4yvIONq/K3tXNJrR7tZQgqY6fVb
u/3LT4K+S7EzptN7Yd0KngGui0KBkKO4o9+Hn1cGAei5OP/p8XKBxkFEc5PE
cwW3JdvonmTEX3AvXOY5JrA3va3Ltn7j7WGkZsadCmYARuJEMwMJDbYkEY6r
i0kprKDprXkyfQbDVlPpM1b3egVlz9v+rMwcBFE87BR4rpJWdqsg4XbqXaqj
qHVYqrDcuMPVseY0N18uJF3OzzSxdzcL0/pfg/My+3w+noJFA3bsuc9c1Xqk
+DGqXV8DNnm11Ov48Yo0hcJsILNs3fkjvJmBWV1AaFmy8Rw/8g22AvYa+c7Z
Ecp90qs4U5BiWkV3vdilHqlQZsOGKnkfDiFgY1+leKkIa+MfnX6RNfswEEpT
sbXCC2t0GJEUr4HZi1WW91TjuLQK2e6niDY8W8Eje5Q02+vUJoYgo7iu6lrE
xaikbcZhMWeIQP958Li/zxJ+EXK8QWoo1uHGJ5nlFOjGw3KiI0vGUWf4HIrj
az7gtoOq30R4CN6Vr5M3B6wFxeZRfv6HGkKSQ/4K6kcBEPvlevzh2Bl7KG+Z
5wDEzsyLfhJd2g3FMaCwyULbtQYEKghLXflmje4CMeU810OAT25hsmFCZ4pW
OQucaDsOYL4T4EWo9pMzbDxzkZQjdDZq0gHaQX7YLvjzzyFgW/dR3sgJiVwf
9qyUBDaJd/N2YvTgNSDTG1wXkNdV/xCr4Hu9SS5Nk0jPnTxspwLcBwGXmdbJ
4F2upPxW5X0ZTNZFagaxvFp3axxzxx40tuP8BBRaoocNMjxFLG4Qv/sHZkfU
wKgMkLLNHf1Z1LwjDO9KFAubGJwfKWmDH42Ok2pAkU2tUpaNBaydjbF96wfb
BC3e1GVRebdZ+MgEVPB1mg0OCi0/+oC7HCc6K2Dc0EyYC8Yl/isX2cqhe3Gg
k4T4I7Gp6h0da4eD+ucEM1oQyfLNefq8rRSMJwK8vP9WNIRN30Fk8AQb2Hqf
QXU09Dr93Dko8AAUXsGjhdCowfGTuQcqU2UsWNk8hc2wrHxfq+BL4Ac/0VQE
zK0X5eYGJByyTE/78ggaEgsjCoQBgudQMtEozwy/uJqX9RlWKDLyZ1mBD17I
WEhEOJcOr+7/3C3LCEC1MsyOGhOMSw9yisq23shshmjQtXI0ky6mJYSEkcdd
X4oneooV/CDOYtVqKzxA3KDOPqYe555SpjtsQn6ZUy7LqiIb8QwTxlVSLxn3
JklY0n515mnFLfyUeGS/NeKyvYa/VqujHyB7i3m8/2U0u/c/mL3Xd5HmEyrw
nUPBefqD8kAP77koYfhxWwL1uTyHvpPnFGERd20togMvVjlH0YsarILTJzcC
9Pey6bJv6CvdqE0o5ANFREUfTq6LxuFbmPjnWwRwUd0JB5XIGLdTDpSarOTW
uWXFZBFVvFN16XXjBdBZVV9Bl6ZI38Zi6Lh+c73d5m5Wg08LGFfxVCWBGM4X
QG4/npeww7wLZHOFnKY8h//YuqEXxqBJnx67rghV2YQFfJpO/GK9sT1ztqmB
7VY78kVhrCHHsLt7GX90dlSnZkBi6+txIGzJsNvR2MU2R3X58ntt78vGSXyp
4z2OVhKESIh0Y8qPEKSF+OgihKgNgeNNxVXoDFE5jvzsdRJ11Ul5YSB6qO4j
bsABd792j4yRXIuDovwgVybnibME7aNrOcUzmMmu3lex1zuJxfCsrECwv5tF
WWHvoz0yqKnOf4AceYfb5VanF0Gf7oULLMTarMTQ9BOONANB0W2lRdck6j2p
4lO9QD8Y/aF9djFXY9QHnlbY0bsnh6j85xSTgEpAPoggMUrYK2MTDcUhXARG
8oTZGj0ndM3hAoiS3TNABwTOPulrU9kRX4HqejiYUXHThFee7/4B2/QQgumz
/kSh5n0mmwMRDH7tdEwrbMWxslIpOzpSnk+KcWbwCQax+8iRJExBGhQRB39/
G4WBHate0+Il/A3ivxfvrG5qX0VHyYM5E8ordVRweBMU9Lte3yT1aB07ilQZ
k+fyEvtPDKyp8jBL0cZ/MIJEDyZ24lm3hbBXO4vH53Akgj+Fu1D9gJ7KcvZN
iX/n+xoukM4I5T/Ca9XAL6cI+bwkB66boB+TA32Wqhasz/OhBST6RhFeNhmf
Mim9mTiTIHSYg+tjqVKsxr3RsFqLnMoZjP9jh35I5e5oCfF6DScLa7glDztk
kR+RZhRA69qOzPoWM5vz/HlwtzV/xqxSQ7N/4Fz3/QiiCjbvfxb9e81uw7x0
dJxY0sg9qmdn4oobduZBRuB8nHu5aYFWLSL4a1Q13n0Dao4tsZQI6KPIX5yH
F4QsXz4L0wSjawqDoiW8cvLIEzZnE/7Kv/CVLzHCepY0Mz+bUaarEnyLQ66A
Car/lwkcOGpI5T9L+SDGyzWhp5/MTpGf9L2ZYPPdJGMur+Od6QkVqrQN/wjQ
wr0mmdisS+kPMxoIJxMejRQWmS6FpJJHZW3xHIhyrB2zH+vFhUSt5hnIC76h
5xkIYzwGkv/bmutzc7IeEj5P/hGoPBK7LJiqIcadOnRuopOHXmRfT8QVJc17
4zJQjcdQ5lcKxk8/IKb6O21wlatGWJ9+5uoG9tEfr014ZcAGtMlrKpDAm5nu
RMrWWGZACjbjtdP/H1v1XXjKIs7KBTXE/1xmpLHuWANaeXTdf9qNIxC28uq0
GCKk1EIzdYnQOcL+4WuVGzV57Cx2DHFAw6JYLVmNZcE7zfZDKDyuRITz4AM+
j1vqbml3Ud+bowpKe3Hf1y58BfEilj+197Cq7DtCsEPNC3Rzn94LwwQBVCQy
qpmMB7rhk95BSnrj4l+wFutn8FFFun+8OZda7qLKEACDsLme+ihK6LHBFGbN
1WOgP+629oFa48/iYlU8Fn+uQxMyimO02x3Xkr6O607onlJuQNaDDMo6CoNY
/wPTmAZKcbDsYBJ29d6QZpy0Tj5pAGFiy4WFmtVOReP7BHbunYq76BKwrHVh
YhRKtJIUf1KnEzTg20nGC1ubk6K4vwAsN+5Oy3CcEsBrGh//86rxhzK7ql28
YwXhZbaa5/jT7VAe5PcwkIqcQW42tUBwsgUDimN/+cwx0nvt79caBAtGo+CZ
PC7OmHHhIO/Qa5kRMysMkSPFlJ9JXMLHUuUMA06DZgM2m1v2+OjeHdxNnm76
1c3HYDN3xJR8HtX5w2pLbJFQKIjke3f1VHzTnDLQXQMQuWrPKLqhx3LeneXo
9qw/xDh14mxlm1CRSLkGNirxh2pGxQKJXYYMW+M5nGSdLTCAh0JuqyEo25Dg
19EFJ3OyLxP6e65aPoNuOFs/d9DfT17VCHt9yhNRG8cuLEDcyoOkJapLBM5Z
k768hgRzXZHaCGGQo4OfEJK7MffMXpnOj16x5qIGFKMr1CIXfqRUus4BjCj3
3wonjoYPd3mu2Ju3tt8nsK1yvCF0i9hB8Df50j4SP/5zps3T/qmJB/6Ysj3j
+Cw/1Mg+4wkNnC7aJ+LIjZ64vJFNrhiIkQaXh3ExRLkzNwACkIS0+Hfmo7JU
QiyimIr0WpI1SVZ3FHVUmm7/j5Fy8RsqBiURlCAz9lvXdgzssQJeYRTyyLgJ
ENiegd9WCOAkkP2zBnME9BTT7F7tgOVkpu5WQsrbQ4kRHyF7Uhmi3D6pSlnt
OUg+2AZSjA3vTFoWEeodGB4arE8NQ7eEaIDS0gBUtbsTKVWj0e4j4ioE4Kks
YpTHRgGj9kpJEbCwe1kvrxs1jARkgAoa4jcwAo4FYK6fP5/kVl8g5kxlJjDo
4kzhgUl1vHu8ohLWG0T1McR0GaJWifQs82wRK7wlujfM5QaTbUcaopOZ6aY0
ppVWurIa++n7bwl1e7/ZATV70mU/pSHyGklX3kSpujraAx+RurGohRMI4qY1
pEVbrXYYGpXaLbBKZB5ld9kA7IBoe+EvJIL+LIbw4WFgwd3iJWhrHra2adTR
QzY3rgmpBdJ5Y39yv64BKaPg1wkFxuBPy+/DMexACSHx03VzeOJoiXFHCUFw
e21rSLq+Y1c9O5sGsYKitZf/J+F3x5mIptoU0sCOkK2ZHuqarSTjnPOASPi+
IrYAIzlek5Y7eKmARdeXQ07YbUiJvyzvWnjFSJY/Eu9xI4ipYvEZhtt5gxHF
xNt02her+StPokEAQBmDl94KrNGCSEw76J4Wbw+JvIUiUOOlFW2TzGE7hiyA
LigOB7EclES1pPVu7neeq7bkIsICGYXYc3csdSkR3XULm7XIklMm4v9HEGNO
5/iQU/YHHdQ2e4G/WE7O8huhYAXUXD/2XczVr2ePZYLp07LJG07h46YaFiTG
CChDemgK/ac/Vj7apPwbipWHaoRIgXjxoAGkWteWsYw23AittX9SfB2GlhqJ
FbE85Ag1Ibj888npD4eeDLOImg+N+Y5pLfrOMv3y8VV8DygyKIkPqWJ0LDIi
d0m+pM1XLyaH+387ce7hjcClO8+JbjkLonNAtU+Op//I+Nb7wEfe80QUakRi
92RXG62s+nsanNhmwlvWXst8W0I6pSdbrVTlBq5tYlTwuuXnV2GA/YjAHmby
gF6T0jUZB8Gdie2RRBco+qB6RJx0AzySecytLvlQwKmSy++8aeu18iefIcR0
z80Giz9hLinI6F5F9cHooxK3JQdS5f6w1Z1q3wBn6bbnrlr2UVpibQbRRs8e
J9f3wLSGKMDuyH5BksBI8kNyXOVbbYsKcwIGWfo/onIK7UWF1TrzmV+fD36Y
BcHJYjG/8TVTtJoWARnjjFANIpHVnHeg2FiSBY+3ADeXPJGma76DChKJVCgj
4r+LDQY83Nb+6ktPiDbsShjF+N6vzDRNMFOZnfQrRT0mbHqYhzmIZoDcPb+G
S7HN/NQlnRc/+KmYlKJxxMOhQE0jApS9uZlC+1m0IFPNrgNOYD28DR00yn0m
1CM/fZM9ISyheNBLqqK5/eoAnOAT3aaHFTQIduHr+lRRsrTv2YMWvnyJuozn
0jGYfbSrzaBXW1p5v84bNUit9h8tjeYyvGw/gf6apxBNZGtwzkZ0qnYHn4TH
oiPX/tpne1JKaiUvjJc0N9LNgiMqWKEGDC4nXZlHZiMB/F17y0KKIpEsa/sg
Y6KjSYNKKRLWBgPlIYYcQnlwQYfSX6wCIPriWKIqzw2yxncxj5OIsLaqhEyb
oCg/v4jB4fD1QUxdz1q86oiaNkQbDpVkBpriCrtm01QLULSUw0fewsNok3jC
FEBVI+CAQqP8IXL+GPRM354u9CFCqlDso7ehHwhAa0Iu3AUr457VvDCx33VD
5VqyMsoIek+meZz6uppXJ6dtTyuLq0KjK0uqa6mmLllUDdIfdznNKODQh8/U
wWlAWKEF2NeRVl91oNw6RKk68OpZVMRMSRY3379n4m9FUiSFFvk+zWMtv7KH
2UqpKjvPKgPUCiMGEWIZZ1Z7gClqbDu8xI7wKXlGy4IvntqkeYjhbtRn/uTw
/Z35nSvwqnyv1mweAsMOqjcljKZ2RDHSAKJeRQfK7lFy/NqXUPbSf9jk6KIV
D6hTYM5L6TS2GTIGnLhEKiXv4bQJCns51J/hWSnbS08VTGSl0mDiSGnnqmO/
u8uQsdYKs+y+hyrNJ37xqhlnr3mEvzKk9ulhbSi2RhCUMfcwmbKCqkLpplns
L3jnS04fXlJMWym0/ptGifFrAS2J71VjyxFljemM7ymBclt3CXnC9TAKNw2o
BpxKtx+AtpB9WMXzaOHX4p0oEKk4gH3cooxRzyPOwIVVHpLEH/+wxY+gbZO+
bzZZeMg6eZ3lbQZTige+pPAJy7lsBkpZwpetmHekxFYS6Kq8/sEMhfgxdXPt
Q4jTG+qJBXq9fpO8ILN6SWjGZY3dm5QX7acPBTrb0iH3cmjOEPUqjFIB9tlq
wZxwVl/aYVVV7ceMtCNbJ/ARJ+bG8GXPo0Pa1MrWHZ2ffxzKduLfZ5r7Uhnx
U6o0cMIVYOihnNgEGv07PleWr51SOeq/bPeSKnJwO6oVy2cY3MekK6qgc+k1
cOUD4bgkFDKUtoxJ9cDiDBm9WN7KUW+AiYYMJVrpEcdG9KwkwIih9W9XCrtQ
d+rXOlWzhFf9GRHbDNNeehBH64tTY4IGAudqxkhFizEqUFMdL0jfI9egAhm5
mAKry5w/kAQcfq2g8Bc2K2T37tUB44r3d8YREe/LuL5VUDmXxBP57ArB2gvj
mlsNeCogUimN8+YNTuYZ7mOtgxxq1oMDTNVGkId/HchaZNxyFVE4N854twxA
+tzfyg55ZwhLX6WDp76AIhbWZTp9tD8MDJsvyij1ifDPFYHiZFqxk3QB/4sh
MmeJV4xMdlgI0rUSAfl3nyA1Y9Wb0gyCOwsEYyzgjbQImDLu9WBGaPka0ElP
cCt8psAzONqZQ5wdmqYSi3SyW5SM1NzFpiaCbnp/oV/yWh63zojs+TZfpUUu
uqHN1qhv4apgA1vshnPvKFjfqvecmDmIP/cZxXYZ6OWWMIt6U/Z+UUZGMsYD
iJ4wI0dGY0S8a6LtHO70NahNf5HdgJ9obdGzORtu5WOcANJgAL8ysu02qDy0
edLQxUy4QDTDCI8+gyLQzwTaZ2JZGWiy6sQNQvwCkyJGzSJ2xJjb3sG9GOk/
4LqdJcKOvuIYl/bPxMDxL8S6iDGBl8h3GDYQvOrexBCQ2UPIbHhD7sOWleYJ
nFHQa+gpnbEPA3Bp0h6qC5tja+lf9E9HChg69E4fUniw2POH9dVbIr4DqMgr
naxAe+VHfWGSSdOoKKj/dk05G1Rz6GmZaLgnxW07jdQSeEIuyS0yOyoyHOjM
Ik54MMk9jaj+eEIhKW7hzzFM0jA3UHn8z/TjJIBQhlnxIAF95W5qp+wwWj4f
At6hIE6m3e502M/Fu/8MtTiKboRbdJiAhm3pGU3gWxVJMdnfAab2CrFA42/z
mljz+3W8KK7aeuqlN0oWDGvguUU/S4FyyjPYpwV/5j5wsbxpHEjxiriiogaK
0pV2WQRGMHTSqXGvYYEdAOFBn8Z1YjofJF9JFGQOFfU6lur0/TRBwEtWUjeo
Wc6M5dJN5NboIPfPnuEjqTSp1USWYIZtck3ANoxxUosfQliEzFCmSPu/MaAL
5N8rpqzMfZCHKBsSr2XVU9AA1MpLiSFeBgl4xJ+MVEeM2QQb2dJrXVEwNhe8
a2OZvR0+yqCL5D1Xkjz1B4EUyjf9m1EEZUpgYfe/nmZormi/chHcQQXxahoM
lnJ9bJITcDML+1c/sG2VIWuzA0ia3b+nkDh/bjO9Sp1C7GMW2nkR4cxIrMeV
LWgLLRR/7EQ2UbpBMD8/7W8JuTyHXhS6WEkzTsTEBbOC2fZgvPJpFWbOGomr
UyyrIQtFL4LIVt+UUnamz/a2R0d1d1G1JOJqaoRE8qep/vxInGBusvl0efrt
wuVlcdOf5pBs+0pII/VViiNww7jPUo7xnb2nh8L/OQgNL0xoQPKHxvrt57AP
RQHUO5FjPnT4yCSgbG5PbOKvrhL7dYrsQjwGk44NNnvUycmo7y1uhc6r9TGs
PFxOXPU6yfO8GeJ2L+mnjP8oAMqBM1y4urOOFpw+1cdlKnOO4VJqYLMEcQ4F
HrgJGtKWVkYMxUaaGkDj7Rj0kga6AGrtLmiSjG4845WxLE0AYHUsQB7bFcCK
+1Bhb/ZL2WU01EelITY7lK0k4AuuNIVjqJ/om69JJYkN93l4MwDkeS9Dr7wd
Rkd/LBfSbyL6LGhE8+CEWSG2CXeuGMCA9Q0EeB5b2dL/XSQmqUk9SQL881KN
Ce5cJZd8vflxL0tX2QX1bOTxB4IKtpB5XGZyHvvfuV78ijrNpd3IgXA9Lt98
Y4DiJ1Z9X+TkzJmn2Oii8Rt8Qh+x4X2883TkMmpGdjkXPbo5xQ8MzXxp4rYJ
79surghkoADrQs+1hBRkWyQa8iNY6aZawrGjctm+JJW8memVzVsc9nIkF5jW
fcsa2gSQbWwoQOIQxaF6wfr2/QjN6UnUWPKQB/Xu/7w8nIbvn4cccbS4UvqV
Mi9OTruroSTcKDvd0BDvG9lg7v42XcBLZ978lwUdrZNhDtSQm/64edGKLsHd
QHms/Qb9nYcw4W3N6WhYgArzD6qNVTy3tRVErYSU4o5Jx2n5vMyq/aMrGGlg
OkvW8+RwK/gwtBj+44yPILoMcOOUOBLa4iCEhz5Nr1nmtLcWJB4oO4/+JWIF
XwwJOT65ZqHHd+iyKswDQT81n735sTBMuh5IN2vViAT9XjuiSzwgFnR/sWxQ
STiTnab2ikbXv3iToH875MdsEQWHExFd0UBsEyQV5oqGBDprzmvJPiJRKjSp
SGf9OQLlXlFzUGrz471NP9nQeeg9MHiTpKkpgVqeVTxU0rZY3Z04YLKgm2nM
XFwxyrvQZfJ+Cfb7iwbuSo/ZVX3P6VeTzUZwZuXe7WOAojoeuRjqrjbxHr3k
QHtxtZ1OtoREEeegvkQntXlyuunw3wV2PTyUQuvZ+/F6awldBthuaZjpd8Fp
5POMDkTXlzCCrHwP3FYewG85/TUnNTB76UU9DuLBEoRefo+ZatrnGBtD/oRU
QpPAWzdv4Bf0cZLNJO7o3NAMhTbn2k0wVobmgJYt10lsSaPuhsI+0aQmHwCf
hTYtqhGZLZw+7ZVvUrVANPnOEfOvIoxT3n8HarB1eXG/+Oc/3BA12xJ8Kl2J
WybUCMvKJ/nk1PvIZyk4pbc+BROzGX1nX8+lePnSDENSlaLPfZih+Na/qksT
4rZDjfQnl/dc1B0Sh6yZlKSd1LM4rfMcGyRhCCeO5WiN7Si3LE31D4ReuEpr
EoeEIc7ppEGUIsjjJNhWp/Ng9CtW/ItCsZldZ/R2RlzXpF7WAqOVqkf5KgtB
oV5KtULKZ74KA9scaIAxQJ9eBM14Vbcxoj68RE4sIdlQouHI4lQSnwRaX+xo
ArFq9ZkogN9n+CE6+XNt+rAISp7TUIoBkqc7KaF/4a7bgSYuHtiPza2v/SDM
9CBuXNTLKEhCf8xAwJdVkYAem4ztXUDX2w4Dy3ZgGTEzZ1ViQT9xQOtmpvMg
fx1Z74JHu8+i2a0+DUZJeXcbeF6HVrwcU7CohiEyZqpQzV3y9a8rC8btG/TI
osl7tk5Dxhyf6KF9v1lCpxnQIh10qj4BQiwsTTlF6WlI8rWDRp4TchlqOkAZ
C6NhuEdIEafjxrP9OxpRVs/+8cWkJ2+OUXsAlDBxg3c91Jwni5jePvmq2Xl0
xKDFKy59dX26pJXeNqg1NNtGCRRHKqlwvnGJkPGWV/qcW2LzUBEtHck+05tL
hwRG0QjmQfqVRzJG4RoktrugX4VItzyPWRbnUQsl31tjTVtrs5KAL2PStyLq
XWS20N63QWuhjU5S0MezKGaCshk2tm6WHTLi8QcZoAb1YpvgEkCtF1r8O9EA
4QC28HdJ0Evj5pmLMq1P16U9uiI+joKZwjZChWC5m3Bl8zoSCL3dabypcE56
sYc0wiIYctnKvq6oUfpDy94ZiXWbieRTlcIEK74aJThrGo0SNm7sfwEMpmFp
p9R7ZV9YOCG1xy8PNq6h+CG6PrRiTFHEsz03kfC3WI1oIU/bAC82Uk8XmdDP
xObQfS2oAeWsMdVZJI4AFiVSkQlo9NfKEWKg5eI/50UIny0jeiAlUYCw2Bhn
wKmgT1Nmfzs4Y5NRVtwM5UOSqegIT7NTSDtaBqrk9k+SP0AaiMmG9XEfRQ+k
Cu8rzbZxZoZVHXMaGC8ohWmCZfFJGVOqHvCodlcbD2NuII5EcsCLEqEEmMFM
/0rL3msAO8+wptKX4dCl4hSbtQPXLGzQG7chPriTeEplRObNLyTJS0aO1W7u
nrx5hF9frGZzkpAvJG7pjb9WpD4vj/h0bNgKSHKzGEKQsN4Oxsuod29Vfo4T
LjKp2IrYd6IacK0JSgw5Kw0OG8N6cTfoy0SdyWOOYTbtNEeI5EpRwm5kRjqA
lCz1/qMAgPmcifI7TadYT5xEdMeaHMoenaTzisU3e5pFfckUCo6M32XsY7ja
w3mYqWCwh7HOg8dwfB+Xw3vV5jmIz0Q1t8FsBpbDDWuQDviJ0firnZfHoVK3
TYtKTFKCDrNAgyaj4oXY7P0MwhAK2tiD9YR3QGFf3EPE8iBLd03GMBl0clrH
UfOMdDkgb/8QrUnLDF4QsQS725IA5+2eosJh4gD6xmxCWzqtwPlzTeU7h8nW
y5Qy5N61UiUG65FMkCQY6j3TiJsWdvQ2iNdnU2JmxUn5NwAXd7dFMLIkNjKi
vJvRsjAxelTXtpi7ehhLnb2oVEk/9wmCSQm50tAuy0XDwSxm9v/6hJEDAHuP
iS81zL6IyhKaI8HnuCTe0vfC7q5FFi56T09miZzIfV6VMW2aBQVEADDBVrZz
cADRAFLOvBQLt4OcomWPe5Q+FhCbgbXlKRw3AGmaXs09mQ7Ktv78iLAr+3Lz
PtA0ECjlhsnkXFepd+MlBmItneEEeGDHtGOzqdh+XVks0LsTaZrmYi1xvHWs
Y53XBiZOTwgIRKzOjITgPC18P9go3hC3Ko5geSlXblOrx5sZ/ncWCH9Xp5hz
UCLAUbSURU9MSU0p/TPhsBZskU75b6HfVoPBrtHCZpTPLfKmKVI5+d2Qvl4F
lBv0m4byEZR+XdmVlvQxDartQJeQwGqkLErE5VM9U09s4uIoroYEvtIguHge
csu8zT8jHycWm98Qo/eBNeK4LIo+gAm3IeS0ivgwWmbRuwGBZYygp11OGU0/
xDQuK9Pcn/VBuPTmzLCOovoLFV1skm1z2yQy/tqv8Da0dteewSXpThYYYWkP
gMvQvjEXZ6Mjl/Q1lPlSMlLaqi5w+YdFmyKOZ5Ur+qO3Ipe3+DFWJbi+Tabn
M1Z+Z5COF3G7a1oUFh+fsC8bMbFm2P7PcbAtpX93YbBy2ZTPKoSY6dUG1Ytu
TqNKGZ3dUaqs9R4SiP1BIqLAs+u7jVFCR/I4BnDarZvvL0g6N1h11m1F3QJU
9lwXBAVnhRCCsH8CdeKAwFFH0hj0sPxOI7vg/8vCJPwvNN7C3WJwBzMJmojx
V1uWUv+vLugyVsNL7bzjJRwvzIxqSH5L7C9wEanReODXD3YMkAImRJybVnaa
ivadIyn3CPgojwLVi0afJY3G3QIaqZHM06VsGynJDz+hbqU7cV3GenUHjviY
LfjgBbGaLkNAs7fzQ4I0d5U2jykKuF9eKCsXIs3N5J7a//waHhh1GrJWsW6c
sJXClCPOyXmO7eq0nCIAsVafJ8YBtigLIES0a+awV4wCeCOPOs7sfEVzrzXS
UXeSRc4dVp520tNUY3X+g6ln7H1LqNLZnLFyCRTmE1wvILAjESZC0RW8eiii
ofDV0oMP9XMXiJNoX9XdORd/tIEJL8aZAzval0h/Y0Ck6FwGDoQqsBiVCa/9
4g+ckRs0/HIYB46KN8uonaIgngCoR/UBiNk6zRRdXYHZWp/PXWMWiAl6Tf8a
virBjNR7X3b87t6jMNb4TvVkQAAWCuch7m4xTQzGl80jtUCrpuPDyLqO0lGt
vqG6Oyfh/NtuuNfY12vMZWqIJDQ6vRbMMRbHYUTPTyBvTxFUJk/Ftg6OTJsj
7Zu2eYzJLd/PADIDA1u8UCWrJbAvXhcF+fPTqd/vyBjB1d3BK5veUZ+8KnHl
xyGB6sUpFM1SBpoBZ2XQtZmvi4ZBibb2LJdP820IxQ911CuyjLiX3nPo35rA
eR5rXmvhJVAer3daY4g4K9/0UymzEQ+3WG5Hq1dOrmNFXoYvoiLgOwy2U1kD
cqIHt4bDGornPjn9zfhiwvcM4O0/5UPz2YG9dsaazm+pIE5oRQNFVnvlnGaj
XpEYhNXARk/oQH1YwqJpqRdvkl2nN43Ql/tryk5tBViISf6rSzoGbePZufiY
U/6B11O0vQmyQVeEzncfvkVja5l16b0P9dWGHUldm969geIR9LAadd+CkEsq
oAZVKmSTsVmag6s1gg5m/vJfHWO4yS/24j8viLc+jeusyHFhqVISC8aWvat0
VNEZ4lBnNTRlORumt8LM3PMh7gTCnT1X6gkQE+C0JvdCqnCxbI4fmwSA4UwX
/Yozu/9PeHyiaxwu0WmHHbCckgm8pSzEuXHOAQTSS4ud9alx4nDwEokdUd/x
Jcepm8LwjE3As5jXVBQ+PClju/94fhBxGq73q+3XkM3OF5+5OwsNA/XCZDI7
HCpH6xcPrwQPJDyhhbSMu/aAIISogoiZ/gtdnFAVmKoHFhgRRfkjbfzGegW8
sMr6VoR9xXwRLp9fTxt7aYraUdNJKgwMlTnFLxswUYDvUV57gc8ux0njm7Q4
xH4uaTypScCU09ThJxx3j/9/97eFs+/1IPpnJ2OoY1lf41qm006Sp7ELniXY
7MSGSaZ/gQ5BGlIXYoAsAiKv1Vp1xC1w8RgCQINC/BZz1a4vfkQQ5XY6hTQI
0T6MY9Ql6h6PXoBz+bWPjmXaNgSvL19AB1cm2cuf8uYZDcbSbsODkWctxGXl
FUADsIVWwihJm8ApQ5ftlIXWX056gNuG2AUl7uRhtjYtZDEGBfbawKDeviS+
A+cqHiFl6h1Kg8eG3TAkon1hjG4uynUFvGP8n1YGYm5lCpW6tdq6JT+e+/Gs
aRi2JlQrw9a6e4q6WizLznFj84Sb7NTMaUTwfV/S8Rd7XFC4slrSVW2wR3Vt
rRwFhgzOPKRTg+HYs2Di/91/9lALMI+SfxeBfNI8Klmy+7iuB+TcmSRz/T9a
OhbvxZtGmqbM4Vcam6bhEWcFsbhrzbei3k+AfoAfggIhYnjZGWrAjMM2ngbl
wni8W7MI4ETVoG4JnxhgfdJQh1JpPyaxV+Z+Z+9B8gnixzLuNDa1HvWKIqik
YTRdiTsMAeCuuNpOiwAyCSyL+FLh16njPn6OZkRdmVXoobgTtmqua01Aq3c5
amLviPAvjfb6ePiRHSWs6+Y1/iXVe07I5DOvgPIVq5/eeUYMpJ/Ibp5Kuh7m
OMVBKXzqiGLA3FwsCIbgT3yHtsv4h85y9avvWaKl8mIel6oH91gG971nZlS2
CMixTHsSazu9zbdwC0UCibreCKzWvCWf8BkaRk22sAPcLnmE7WqZOwaiqDJ4
2Cvs0UtH1u3Rtw9SzxPU95rnYLQ1dgaq7Y2Bb7WYemPpEOCL9dWwbQYiR12x
R1sSERSwCPSRa74orA3waaT0qLFmjs3T4l9cIUQR9N8D71A9I4mWIqeK7bZU
wO+5f1zUoxmBg4nQvg73j0U2UdAlxw7GLwkJ6JBWoLENPhxRj4a+o3219CNi
m59VnQ8kksMliyZ8Z0/G9Ust7GvM0MurT7ON1R3HkHCUZhQLmXDnMRtMXFQK
MWz3b+CSxKQUjXWK/lN+A4HX/SF89TLSnKnybxftLLReUSg5muD3aSE3/Hum
suK+/t1mYarvDqeA09uOnHRtbRp2JdARCPX2Kvf5PapBfLUysj80jG3HGT5t
4VdU8BZizWgbMj25J3Sp/FcMpR8/4GPMPSXg63hkZAzZvAhaLvj3kIYIWVVd
GC30UN9iU/K+waPlP3Vz3nskudJR9rfvhs9vc8ndZrGOKcdv5N1H+YBtIcq9
mwpmcybP5A4aU5fcKVoPKU3AhXhuqvPdKK+0z54actdzJvgxZSxuG6+wX82R
oA9Pc9SmJG9Od3IdiBrTUo9Ad94toR55Xx7lzQ/6SYQRZDoQ4Wts/R5XKuVH
mXTFeznALMDmP/pgw56HOsrtYynbitBBo1xRPSywx0IZMLesncrQFJPKHjrT
qmnj2SmVekF1xZFbYsGWH4egkAIQw2flIRs04dSOd70TQulAW7lfK8G938Dc
D64nHCC+DuuwOlSLOV3Vm+NASUFumNRxeq92e1g2kIa2FUNB2LmaOhgo8top
MgJxF+57KkYw9hMF5FtoXbb/B3GxLLb+IPrEgY7uCPrmnElUpSYthSQ71B3/
F94WdAYb59JMhNHby4GO18ZcKI4GEg4M9ujSTzZlv4ttUKGDcfGXVYtVPKoY
wFDHcCIVsRgVUq18hEfvvN3ylmee2GmzbyJ+Irj1c558zWTyjVHjKkyFqumE
gAUAtOGcCheVYZ5V6KrGs9TG2YjfrrIGsx+kwTOKRMbQLqrESf66xL30k5cH
f4QPUGxZriMRN6Yqc1fhnlmV2O+pXsBwY4FM74RpLlb+ogeiVAAb4EizCa1G
kwvIbQLM4aitCnH5BLwlR+xFYUHNp7eLK297ElH0+514VDTFmpDN9peSywkO
hwVwPv5IW1nS6heg9Lg8XKVJn9b8VsTfegyPpT5wJTS6AMYHoDVxzU3gZ8tE
msX+k+tqkggTZLd/Wh0DP2ikRnSWDyc6MUjyUDWnBS8nd7x1/ivsqB1F8EYU
WyWvPJBZ7hK0itYvlxIt3bxUtQ+QAZ+4fcknVdi6lIPSeZhPymk/s7+X75HD
Uyx5GHOjIr05f0rhJgNwKxpefomcSJjl93C44M6oF3PytEaU4W0NjIDkTQEz
gKUG8N2BQA6qTfT0VsskVBhhVG15apPTRJZAk6iPQAzlIKaQi50l1WmQA95z
eBdfk7rqoD077u6sZwLpfg+bVQI23Rq/bB8aLNttk3xaBM1sR+6+HF1d5kvo
/BmM5D1/IeHSG7njKhmzH+4Uu4O+Dyl1rMEiJsBPKCbfRBhdgbiZN7/eozJ/
bxb+91sEDzw8MskD7Swr3/VZSWjExgUB8D+K3QqIWD4TZq4XeTnxc/k+Nn9L
42Tj1XhyRVgqzaswo65Wyqd/U6U9HiC8jE7GVm3eW5MGGUuRem7Y/vFisomo
I/O7otWThAYvkKM+owyV/cIJCSfppKqeXukrYW8daGwNy+0/SX59SOI7Uk59
Gi4TtQXZy42BI1pPefZJbzGzs9mviTGNnmklQaFX9nmlU9lw2PmeS5Y7Kr4n
kc8E2p05GmLU65EOB8MlMTSfmpPsI16J9hACajY+uZAmkdyRNqS78oju7tjF
I6biNicIJtGUIaHzpn1amw+UnjqSYUsgBDF3fWO/ni54nG4GrhTbaoYQEFeH
tbducz2aOL2LrND6PHlshkyvDyQp5dXlOsblh8rjsbak2GrK4HJArH4H13o3
jqTlEnKAxwGNmK2Gx+K1X/RRcr55YU1XAtTXW/HjBbtpHcnI202+cneI4JxI
p4qBEAj1v/o0VSuqbQZaCG2/TR4QVPu7ENOY7sWRFoX6f1pl8bk78M3UfaX6
qt5NnC3qVQOV7FVbDTOLOXp8VTZMUxKB5/sQsD1NyipGaHXLSZG70pe+le54
38QF6giywWn5KAqTQXnAlYtVTSXUMy2EGAdwb08gFeUqudCDxCzprahNUuin
bZuu6aqgXEoETexJ7JY4FziE0JRh6EwHTbsYWUJGZeb8QX0mUzUc3Wv1JJIN
jGv5I/tuKFs5l+C96mO1fF5/KawqxKJGN7oaXJaVmuY84gIWkL/8qPfwVVbG
T1pFDJnp7YrVXe61GGEsMT4IEhcT7M5PlnEMJIV1VrPYmq4BDOdwsdcpdHM3
UkgDlxcOVK+Byy7U+S+BuMCyuD+Eb9fug4xnPeK0hE85bPXlyxl4qWl0HisN
HOsqVtnehaMSHukI5ou/wnkPa/8oI6h7KG4HKmk4EXRgk8TZOMsjIedjuK+B
cR2W+AMyDr1lcVagLShDlh2SGUO3lMPv42d+cSyQ0Ql9xnr+HH3Yqj7eCgSL
ymMXjK0QuQFMheZxX+7YynJjRQDV1yujLneThtyPIVo3Wa/m2Fl58RzQ034a
MER49DN6zagzlHniBSfKAdU/2Cv0qHS0jBdWm7hVlgCOwn2MdiXcV9GB8J8j
iHoxhEvc0GicUpJt1LHO7I/2Tx4QdQfQ3k+ykJsDykA8cB7mge100qtisOZZ
chXErde5TPU5Q/sDASVgFvJM2dTNciKYz2U9xqzvoRzwV8F2b5NwzZxFST6N
B12AApQB4kscBQtIgP6D8LZPRTwfrHAVmwRxblXPKpWFkEQQE6H+QDLwzWs7
NS4Xrv+Yh6ovYaQ/7CmLalLA4YS2PQqG4zGrH9V/yzLDJ/JT8XtDDNDgafvI
NTgJJDN1pFj/acKsldEM98zOQKNXZNaREm/fuAh1KbuhpLAD+TZQA30j0Ktj
0D9IPrvWTzhK50rLaBaDhoSZ7szCbr4MI7NZnC1mJ6eNGNZhLOVOriZcNb+A
VVfTYA/a29Xdm57/tgGrnFxys950jeU+a7NqHxyaa+iD5ckiRE4ksDXj8LDk
WBVfAlb9sXVRHbEee1WINohUlPCH+9EPhaeiuhGn20aS0ultQ2+95M6Rj04Q
2n3P884h53PCSMRmdXDwb9dQUpg1IWFwfZVgxTbvRm3VYPk9rfmo0UE1pK1d
eAZnga63aQjER5yZu8GSYN5KizYZ8rlQ+ZS/fYv01xbqrTc3ON0YKhIIXXwC
k/7/5MK/bH+lc9u65UkSlqk9bRZna7C2ANrZ+BQEh9Dahbi5U/hKdbx2cWIm
64fPQ/fKi6HjCNKZgyVoHiQP3G/1dzWfqUHmrfQtC0kgL3QX/sU33+/7ClVl
iBpbWwyAupsRQ103wdXixWCAbuUjBrY2WgBDPURT4+YT/rQdeIQoP34FFkTZ
G++sHPH01Ul0AuNj5LQoaIfEFEEb5fguNKTTB61K0pyxAMeBvd+6cHY6eQb7
Ik8TrymkoZbHSRiIrJIJZ556X8yJZkr7X50DwE/GdYsGh0diQa0rBz+htTjW
tflr2LnBbhsbmmAS9nO9qEAsW8rkwGS3U0anIwJQk5xCxIAyVmQyubtlD0n9
BrKKJuRNbTej6rVExe9ciuUpmOfj9r9w1f0S7fQ7qYSVDkjXt0jwNrbAEumt
Eio8KpMRD9u762JbzLbdqiaIV1eU+tzTu5jQu8Dfk5iY9oSXl+WilWU2Acqg
JKk0jq2uuQ7nkP4p+w9slFnYQUvo3dRmxT26zPmrrIp3c0kUZr6QEmDs1boz
Z9RVuEMEPIiFIR1q0B8o1PNGuoAIj8kg5OhYt6BwrkDxLK5r0oXUfEFpyexm
O6cKA9fl9LVf2OCmWLsbvJcAsJWfCU7xl6jIm5dnJB+t2NtpLiD8G32yBV3G
5vVSoovhBry7IUtIJviWRl2p0x5/shytqP28Br1ItrY88HH3qMHeqomvRCnL
0/6j+rjpeDATXsDg0WqDYdURfdYqo8OKLbuAgOdtclCU47mx0Moe/78Hbpho
i4p9Z+yAfx1b2S1gDXwnXSY2ednV+1XMlFtUX4HCrh1MTTFOE+qPI8GzXA9A
QBQb8/s30gd72J2A16zmzsauJtm5fpVKqBOZAvxMRliSkEmZlgMM45NvabsV
Wv+F1lP/H1TJRaC7Cv9sJzlyChPW9fqJqTncEfU7JkeqSU1Fjes7HgKWkI4O
zaaHGYybvREoJVyQX3ysBro7mqBTu+1ZGQWlR4hi7V2szmYb/jfTkW9rsujl
mEAbH75SzjwQDarKRQtxF/tNJtfBJYvAis7X5M0TW8THVFrKBEAxAYC6NAR4
vtR6bL0pgcez6vEO0SmFmPTAbZoOk6YtRFH1ynYQFFwCDqdiGbruI6SeiPfP
T7znLpUO6tO2UK9PMYsAD/hw+yEe1nYQNHTr7bLve7reHwTrPlq2LUC8BdMW
rFVme7+mAV6d6kCrxYgAnZ+hNR9SZMnz71GWLCu4sxvBzIWOJguB4cjPkOZL
c6BRR7Rh/kbCa8XdwPd6RkM9SzkCK3nlr+qkVZecQFs7Dw9pulIlXGtDJOBf
jXvgxicnCeJD1AW9Jb9B3Ifv3LWdsi2VaA799evsk6xNF9QVccuCKjA1I+28
QQozOK+XqhBLNM+4N2WQd667qnnoCxrNVeqca+gonuZDJUScfI3/vmUsxV+1
WXqPgAcK6HNE4sm06m6X86DeHRXJcTMJ/LC+ELHGUewgDmBJbNu7fyjZKtqS
0wfRBoz8LI8h8mTBEY2njSTh5uLqOrHiEfw3pO4z9oz+hh7qEAhKc6X8yQAM
DYywhM0bm6yf4BVeCGnouZvGehuweHL+dmdYBHT4Yf6oSG8eJVYkAFmHPrFP
HFfyjsgnpPLITxZJPUIALZsEazyVrpGHGceoMpcoabOb8dwPf/+Wqi9gV35D
Fb8f3F7CTvj/CqDQZQa6ERjyftV5TUywhPFSFCREts7wTebECr7A0uSfBd8V
BxJj9pIx41nVj0wf6F2TYFQiIjzsqAGwaTcO2icAtKRxHvYtyyJMLReqkBX/
e7kHlThxvZ6q5hYobUUMsJnTyz7FejUP6sazkJk+NsOjI+LoZpN52pwoCH0c
mAD1qHtRiNI66WQBdg+LRJBxELHnqrBE2jy6Dw1/F45Ys/jgvvn08JIEd1OD
k8AOpJX2wWNC3yJ8jeWmZZbbHv5WgSlhu+ymp5BEaExu02YmMlA49S1ldTq9
ImOApIN1o3Ze9W8iJxHiH1WfScWt9+r30xHYVnqZzDQMViSt6SQ7OCpyIJbo
LL/I9Q+EmvvlmysX8h0qbhWF4FTEmWjGmDitNaZEbFu1Q1j2WVq5kePLgPTf
X28tx2sWD3x0MzFvNCKLT5TOjhUMZccnWXNFjDyx3EODdF7AIcpUVBFm7eF4
QFL28iuZ2xi+VRsFGvQpLIrelrY/123CRdhOr1NBnR0tLy9mj2TzceQvpVpE
srmqY3+OEJcHM7K5G1XwBkHMFgNwBYIu0hIHmtTw/Y0o1RUsXRF5wovvZIOG
m6RlI4UCu21NxOOjU1cqxmzCC02WKqmIJkyjctbzxbrRCbqtc5z9Spf1KA+N
xrS/Rzd2rdDhsyBRmo+cnqKsq5jkrWeLw1DxJxerUuAftUfIbZX+bO66/oNW
Y1uXtL86xSiWp4bIyDKdzN58995+tGicumw/NlwKwggUQxgqYL+R6wYuMC7E
rslPNwfgYraHBbYNs7Td0E84Ufv9SXS5j2YiWxDmiYS4g2pcyzNkjBXSJNa9
xrNreL4D8OHBlLiNtXh/0Ln4EjSEnQPHj6Quv1v++Nx6OieJPqYeP8K5fGpm
xLwuWNvYCkhqwqru8jnAfTpddUKPURRqVZ94/lMWa2Rbkr3nunNlmu0T0tqd
MJM5eQAW5FOFZL82GBVc9GoiZcO1Y42ui4jwKervXIhqERQ5BFe2RnsPU9wh
V2p5Ijhpm5N4GE86t1dE2GQmVMoeAXlNBmaiuXfC8wWbWPPZTxRwTuv6h2bk
KuN8+FhioDemy+he+b1PowMnpdqKwdOIR2rtBuDumgJyn80dVj6L5wFIZhta
hq2tLKwNpewyWY+03k24sD8VVlsHyvtXtpMAl/gz8onHoeQcMws86ce9ov3H
RI41XEk9A5jwst27WkCtY8rBaEkTnlfn3fUp9c4qtsOPVu/FlqIvNsD8HQXq
VwxvcfsS1zyYSRkUUCier09Sj1B0XIXdIrf+oq1qcWfcTwA/QuI9Km0VaMaz
CxxVUu7FUNIjGJSk8BQyu0NByYjvtOyXHQ4v0JuZqg3CY5rSsOMTrSdhhXwP
2pnluD0N0pxxXYfRnE7deY7WIpnNFT82iWDyudfiIR+yMnuvQqd+Y//jH7ET
E+P/zSWfrdmvbkXoYsItddkhvvhsFbFkEwLb8ZpM5aWie+/3MsaAGYwoQgq+
P71z4agdY/PabYi5pgxYoQRz8+ZySPBLLnQhRtJyjKNFjCEJHl/MowSjvJR6
GO74/kz1pccmt0tUITYhzsuf0v3NIXf2fgoNaNTDcrZg0h8wVwatAAGTtJrm
HXI06/A/O2JZIQoa/F71hf+HimmklCC/Y+2lv/IiGnBcSZNMqt/9pSe0KSqx
I4uTAXmc3RCqhXU8if6e7+avV1rjY9E4VRMr3i1ulRHw0hztX8DOGEYD59xS
rUM7L5J5FWT5V/ibXGjxOndUpQOh1aSBaoCpYefOUlY3A/YspJYXSmUgUvCR
AhMOHJRFikv4tXlyV8ffDQkvnWfsfwdfVw0jl5K34uT93eYIFP77JLQeUZGC
oyXkqjrgEtPINKm/rJvK+ymCDp4S46lNReDsJ1o4HydRXL7KyzSmztEr2oYN
Pu5ZsM5dKeOhnhHmVTrGosnmiso2nKfVYSf77zwpW6sMT4mkkmWzU/aVHALe
nRT/j30mY1n3KEtuRbS4a+rhgab5hdR1rItrF+7a7ELJQ3X8mYdFWs772oRO
k1oID5mrFzKtxGqFVG6I+5pvZ0aygrOCmWb1BIapwB6seCzxWyWw0y6ufrgR
OcE78Q9m95rIQ6z8OAOoMm8NOm6DJxA1ogozVa0X2pQGxORM7hAZWHpUGVmv
f5gOqk+2RddFZivUwWntJLiU4iEgNhkVngKgFSGlhi+1PLX4YWkAbE8J58f3
9P++WJSkV+oA8NDlOTZf//AIKUvwOJ9YoSHdsMAWMsAtYrHmgjVfTKzi03Pp
Vbi3dmBNuC0NPte7nWGKElOQzy9SRRXuQ1wSeNcKBsENNx5MqlxxB2eFba16
L7KKcCUNs7z2IY+HRcNUzGj+6TZVHGZ79Vp4GS6aMh3PLsVNFBi/LQINpBpM
BYqMRk/jxXiUV0hzueJtt9LMyFM1PEikIlrrzhQWaeBP1Vzqvww7WIUNDlMp
bfS2kMjqGZGteBq5OOfkiQnOpXnINdpepTwp+h1pFeFvyvbPko6jagPWuNWb
9c2RgiLkp3W7yQPmEKALHFAkXhqWtkJgE17u17NPwDRKIKm7vj3UdJpWapRz
gVJVjMGVIUGDfLtbU4ztdEm9l1LtBxu7EumfXhrustIP+CQD+bLymc8AEbPw
lfbB9NWDx4yaUa5AAHDIsXv9tWl5PxcFMDhNcWdlHfU+AIkNn4IcOqvTvx1O
QztgkeHpK8sNWNdPQyKN7a4PMORJBfyA8UceZwyWRWVItpsugvN492UGLo3U
KbK9U+Et100lj6QrCKR8rovIXkZc8dYrHi1kW3KV8KUH+s660k4O0UY6q2aA
F6V8pYeW0ZAauKLSXsXGHvMqDfo2dV17HFWV33CSmOKo9jDvRiMKyMJo8YVq
YxHvtVY5VHdkRsXvDCanNfzJMITMiUHi30JSJK5kBkt016tT/+CyJ6xwnNuE
e/dVroozzQd7aqaCbtc5VwJ2hhtFRKQU3M+Oq0ndzBr1IRPcwCj/QaNLkT78
fTZAtUFOkOiyS2K253v33PY9XiPYRDib5mJmU2h+RvbPZs5ZHsvCE6PEnSa6
haRyraggVPZWx5gLAScTJbLAv2JNkLISEepCRPqRhmR3HYE2o5J1Xk3vHWd/
va8BpkX8PQDt4nqgi0RZx8AWlpwgFBw5r1JBujyf7sjVgaFf9ZFH7l8P5a7O
WBhSKwUjVnLDoHDIQMv0zyI55Ps2x1j07gcrc68903hG2AgVi1jQB5sjTfeE
zWrav3/Q2R+NnqLXlM9KnnUsd5bMnp37klHgq3oVyvsyGyvP05MpYjjhRJ/l
CLsOVRDH/rXyID//ejZdJiTpVW7vExalZZrsVstVEEHk/xacPwh/5aptA0iz
zZE+VsA7O0VtJZHA526czW65CyFtJDlH88G8hQKqc721eAavXK7oGVW2FE0L
WFm0Cm8xKM23x8ALyS6lMNrSauoPdavL0MYSSp+5Uyx3r6fx8MRxzZaUwrO9
lS4vFXL/TYO1xLKaCRRwOnIIglbtPH64ow5XuZrI48LHVAa3yoXoMz35zi5/
buVLLjQxKbsmZpqrrDRCwPchydL/uKRAsxAKNpXV8wsESyBz1Uw+R5o3HJml
IbLtV26X2xh5YrNsceFqRgZ5QN2vJGG3s3QiqxKD0LNLVHkWHC1DDnCsXR78
GxWG6ETCYLSGEBsDOigCLLpMaGdDCmW6HxAoqy6jCA/m0e72YXeik65CaR13
Qp0Kg3fBLn+R/tVgEQHF5ahYmOqUN/81zAR4uQj/Y2rBteiTTX0HilBcJEiO
Lw5W40o5aweac8p9NVtPYswfTU5hrAVDRI1MU6EEpv7JHbIWz6h+cveKQvaO
ZmPO5Dx4xYizS6Pg+TKjClEbqp73g6/WrJb9aPnS/oVgE6M1Zlb5Sm965MoF
ggXvU82A2Qbs/VHDrTETUfX391+jkiHzUvm0ReD1BY3uN1SLiohimwWcrKIX
KnA2dWiL/H7KxGQP0HrFxGEWN0x1gBQ46SQpG8Qotha9gPCOHnihNV+bQDoO
Akjr66Ol9NXdDFHgDh8T1kAD/eD+RpWB7JeAf+QufKGQsUErTIuBu6DPgn/o
9kJ39hpHE96sSuEj3fzpeU8Ggb0fUY1MexekgAxLyP6/FsRWBdCvB/rb8eaQ
IH0+IvUHMiUXiz3jL0S/8jJ+vR/Z3egQqdM5rXixKqpa3hoXbt2x474aHmKm
onjhS0xi6NI7mY6QZKrbrXpKkqqVDisTy4DUq9m98cyLWtBfJ6a00A3XTVmb
+LKbU5YpwbHJG6pZwOuNGTsWWuwr/dgZZuNBujyJ/w4o/WW4yYU5JawSMOl8
x/zK35q6mxr9oinabnTQL8aOVYTkf9bSxnZ1Qh/pBG2JIJK0peJ+x4Zks0su
8NJmYDakYWQ0oxWBlsLm/Nvq3JqcsGaONkaFwI+XDn4DWlS/RjNyVO8K5f1l
lC2OsQ2xNWHc7kZT7wqwjrrFu5it0L9vsIqmY92tNvv8sc+mm1dprFfuzHj/
qCXxqZ91cyDvgl2J+m/FuyjWpquGC/m5bpLWRM2Chq4tvXK8+zVb2oKExWkF
cS1FBNCaxJl9uvxPCcL3wPDF+zu5TzkUfOkKJUV5syW8Lx8OwUAl7LMcPWf3
Pe5EKhxaaxf4fbcLD6DWFVwiPL90RMUlPro/n3scuY+TIy0V95u8b6UVP3At
nIFZJ/WtywxyLzjMcEaFNHa0SZO5cQXyQq3xFVA4ySiHHAtktYD9weu88uwp
Dsn2VMq61j/vYTAQsbDgkTLmxR0ssa5KCp0taaCKWKZgVtKKQLHdbHv53cQL
TsqXeJqpo9JNzVFyhLROLt7yIww4JZy4VDFWpU5HDxHMEiuHaCBRJskch0U5
w6BTTo2igunXIY70j++n4SyiLXehdq9ZR7YwzY3xiblkx48C+dFmBLMqD4iL
4vITqwAqSE/9+Xh49korvzj00PDqW8J2NXkLxCYJ3nE2uhpPAGSsw2t1eNXr
0hJa3oYDJRYl6/3BA2ltCrIiQ868zvCMb3nmjbFnDBi3OFd/azhx2H9LcdgP
FPnw0vUAEc4M+dmyGdCDTTOAk/R0f15HteWII0WYzSNm9n8GfTIWPVzzb65O
gu9JDrk8GUMPW1MnPCEl5jV7RwRMLFAnb8DTFo1PkZ8Fcpsxxt0PqyykE27q
ganfBHytJTbLfjq0hEd2j2rSyMcMLAISDVZn5FT9j2+00XcEx0d4vSVmmH9m
4cXNWUDjw/+fXJKgQuOF6vtDo4BtFqsqfCRsFpO+ks2L+tNk9eHeQUemB4w9
BOT1j9ZTzfug5+SL3Xi8TlD3vRvVGojWEe+Ercump2X5kOmamSykZ7nSEitg
NxnZtZe8tzWypKetSn0gk7Erh/v79BaqVjoGt0AJT8c615yOOESRDjoJAJCI
nxZ1sidQ1vF9cKDypND8KuY2Hl4lDb0UCTiyXD6XB+BH4wjr+WPHWKx1HJkm
+LD4/j+nyT7Oedp2yazDV3vsUBgG5F98mogigDtqC/uorvAvZJHIsN91rzAz
EC8IXibt+uE8DlfPN4ff84M5SFwpthzVQLamWJh5IjzSHzxFd6EelVBITem7
wX4OuzTM4L0DAoVFZ/qXL/RTwKoH5isE6HNgfmK3zxQHtwnJk01yHTsNLwCy
d6jQvMcrfu4Oza0degwgqGNz1QFwgW4/OmqVrEnSojO1tQyPfW7CduiIVyt2
yME1dFR/6ZyAIaaR2LgCLjYbuIXIgqi+w9SGr61XazvVW03U+hpfchyUITTA
Q4FnmEwqoeg48Vdhv82LH3sOqQyBr318Y96WpI7ednNMXg3d9byGy0/pCXmP
LuGRjH9fLDR5pbjOi2dXaEZSLFPKYUDuq7FFSBJ4hRxlZNNNFgjGpfHy8Ij0
1oLECYX0nkylbVwPaAf0jKu2AwaJP/urP6ibFMAkRV74I3YT64/Z3l/phNJn
LKy6o8N+80F+3iv5QIAI5GdDokntTHhatc5yX1dxPodP+s/V3MotlDPypJt+
aU5TmNjCwSBdTqkV9TORFECmrmjxWgQ6ngUix0S2FAkJ3IMK3AbPMrisKnI/
b24LFhyiDBPrf/MEgrHRis1vK9KwGqS2h7Yv+3xycDZeokghI+USmsp/vHhf
/07gK8qpUQ96c73NysBravyb4GxwFUXMYFeft/jRuJVCSDY5tdNkn9nOnc/y
YK0ApGffvtEvPteLkXIXt9RenZeE2gKW+O8hqwkmPtPSd+UiDMYgNUkMYifN
9LEIDCTT1mcdzgTNHJFNXqKsTkbKX9MyVJWsXHgWgS1jCBk6VJeiLIyirUDA
23JM1qKIFno9RC5l2+2T2jPJ0NgMURcq78fxcoYrMw/zuad6n3UIzQ42tToM
wBLb5x2kH5wganty2bFM615X3dGiTl5AX23qmr0iwFbbOTsN52PYvqp6h5yD
nM3a3zSFzeHRgkv73JEjeHR5VEeXbNxChP4HT2mEanPPgbVx6ai+Dk5y3+7f
lrmz9EAD5bFohBRPLoA9vr3ALi0f6EYWF/3sLB5m2T29bnR2axyWRNuTsmDv
Qn7zepJhn/uTJod11HFN41Mqtjclpk3fzUWTpsSNZZRMjZ2NORvAavZgEuyf
6YFvrfId6L+q9jdpWswV0vJZmUuZy84syQ06M6o/bAgb8/AkJk+jdTFaieE3
0j31bAuXsoEIoSOsaf3NRSAVCVLU42m1Ow3Zk2u7SBmcDfF7dl5q8iO+1RIV
XeqIF5L6Q1/xi5c5xq9ceGmOLHFyz6Tl0S7DiBkus9XLHgNFXQlI9l2cqU2v
1BcoST0EfMZsCL6SU0lqv9dnNAJRF+2mfUl41grPEF7gE+SFwnxOCyWsmr7v
t8vr1AWmhYPClwjBPaLxue8TcT/jCANVKV/DjVCk0gHEqOx5gm4d6S2eJj1x
rB2LnRoOidaEbkLmiP+4LDaMEUIJ55eaV8D+jTM6aADQuREqelMxAS2ytQr7
Qsg0s1zIeyC+TcBlRC7dKOlMKMqx6l8ejAC8D5/KNjt7/bZaK8kIwWCTWvPQ
OoYH2+xsx7q7PhsXqAMMUZeRs2raTzvj29wK15v4M7xJp6Lu3I+b6bNkgRNq
YuHoNZwEL/CkNbvSG0Erm05LsXjDEFaVQMhCREWcotxObUlfKxoEvdb6KSdP
mEJ56foCneU5G94tT0bw/YXmtnStG2+ig3QfpP7UYF9PBroh6Gn1H0cETeBs
9r5Vj86h4CNW6qKFOr0+K+MIyRW+pg7PerYOA6C7qQ1I6Ox22mzE61yS9RKT
JYUSwj99wukCPGJt2stzOn2JsV0bxTJ/LIiPx0HtZ7/QTD9r6tBqE62uDdHL
xTkzP6B4o6cc8zos6c/hJ2bumTY+8wIsv0UkArjE/U+Ar2W54w7UQY1S8diB
PiXqCvJLAMmz1mQrVD4Rsvh5vzeRPY3qmmzJVllLXjqxWs0m9QuYqQ+LrsdB
H8BEEq9XqVBKYHCwVP9lIfdgE1HwNer9PwFZWAW5zjeggLZgAjeC2v4Q9maN
+9fki9Zk7/rm+J8tTNv7THnqZIK6Qi53S+ijaoDO19AV6NCtDkpCTHz91YN2
/puVGq1TtrK+wXf2IQMMfs1JvIpcP5/CaXpkoR/vCeZKEemhw5v0UArlgzh8
aLtJ121A/KmRWKOnhmHfTbf4BEJ9p/nZmU2aPP+yMMFZyqrPqzHPzWGLY91V
dYfg9o618QmdXEH1jYhVtQ4M4zgso04z4dE4CBZT6Q8LYpgdlnw1Z+oEk9/0
134Al8QM2exRrShRKhncSvJBdyYU8YV143hrIOOHgY8jaV3EzZmw3xbWftk+
D+AJ4JtnT6MsNYqWWY7WKCiDd1ZwASYSHZ00GUDUDvSIIjfZw77OE4qHl9Ic
Y2oX+sdLz6lX6WKHjrxphDgkzd8ZzVVxcfuueGgCX/0Z53w89YVsVGD1X12t
NNu5X9Q0JlmClVIfl2mZqQTuRM+wT/gJYCgLUhw9bhI8GzA1kTbTuTQKkOwq
5wdZCZUXvr49jX9rsNZ03cETuokz1bSZ/1gu07BYBFs07KRsqCHzniqqYLN8
VC8zj+MVbF4J9ynx/Nd6lZOH/Zp2PkJrJ5n2HqvjLOzEDykBhi4iLD9RKimT
shHQRdMdCircUP+4H/rSO58K/j0Btv1sI46FCI4Rhi+tWHfsvyOcKgPzYI5t
jBnAV1neRC/LbdvyJo60h8B66UtQDgLrwWuvnOOMoe66Wp1+TPMUMzPXgY7j
3GuWavuY9uaf5YfSk5lIP9N7uA5Nw+xiss3c/lzyhryE5xmZ45CbiLD0xpYk
jpgK0WB7eflt2ZHJ29sxkPgm2UcRRmUGKrHhvLZ1NpzdIT4oUoe4hq7bhzoU
KMN+PPWL58JbsSNB66WP2ZFgrB3m2A6a5wFwS2MZKFwFwwqRPVy7j7k+yQN/
BEkWFVwy8PoM6hYhwP/12KNOeOygM3qkObtB+nXzWzUhWGZaCrde2H8IPxZ+
UdlInan3aCMHGRZ6j4BgAJ+yha7xfuU/Z2H2i6njj29XjYCMaZRgiSnhzH7i
S15RYhqLZXAfEPY+avl9gOHVqNXzXUTB4zr4eMtnU/uLZTCxMa2JFXnCyfsq
AKSG9ARi0oSiiub8XPOBNorvABh9WmwY01aMxOpLk9k59WuPbqLz79UFdmIA
19fby60IlwR7Z0ICW8MS8eD4wkfRVXOovlal6QPIsC8n98JRnxc27hq3nFAi
zIEKakQEDMA0AOYtKBLN0PyptnD1SMSyJZx6KQIoaZ6+EXthOUq9ojluxDA7
uALOB/i8zbJSrWUfmUspLb6XUwcT6vVzhdUzu5o3gpwW9rzBq5I0HbtRkgWn
F1n1DGXGwWz9lG/UjVe/jF17E7CZtKYNYZWW1ismnCFgBg7N/Ywx1A/SQ+rd
ZhbcJC+3lanUxhe72iHKPGyO0PdPtbI3L5NwHzTfG0a0dZyPq4WRvTrc0HTb
1LeNpg5Qecs6TCrQmz0B9JtZnUV9yU0TRHNyEeGiBsd0w0dMYYkZtBJR91wQ
JH3hH7PJ9g4rLoevzofXOzMlAmijsa2CKCb+OosIxPQ1VeuWxGD8/gSSQaQ7
jhlvf3pAwXyA04jlzveSrxlbJ5HofUoAQurHGPM9/tNYLca7pi2jobWGKb/R
QbjXrSc0nK2HDd0AMky3TbWwPegaYXrXNiMEeFe7fYz9AkY6hp5E4XoSrAzR
srv2Dq+SsqCU62O3vgqrnyhmuVPztUTZQdpE4VblIXmdaVtgsdWj2st+5/j+
K1RHsW/kSeWVXt9rjbFXrrmbv2TDMEL0Gx+hnoicF9qz1uDk00PtpUOk1Xvx
/uJTbLJxMtUbxlz83zed7Vc48jO0DAhI7zrhB3WXY9wCHxvx47rixzsMqK7D
70Umpy7fvKM/La/weEK/2w7Ay0sL7Gg+HHDbBYiCvnpGtmUJjsH6mGRk7hwp
d8pEhBAubgiIgJtSNz8BY2n+fHDLNi6qJXRptBy1y85+osBUNzlMM5RjLXGy
zsGUQ4XQmNaHgcIDu2+U0ikd5FeQvmO2PMK9b4+S6aIkxNaBLi4l6ODxlyBj
CJI3Nt3n1FUGIaa+5Pr2Njj0FLDwzowm+4zjOnVAGqEiQRZSG869Knc7AG6Y
0NFwDJYpHS+SnnIZ1CNGBRbTOEgpkmymosulco1+OP1UiLTY2MM7krL4t9lR
QPPA0TtnyoOv/SPsh8lvNqGypZZreOQWTbLamqHxy/08A03RNVmlYjVFa4f+
vLvgnOsF3ZRtyzcgUwpQ0BPGwTA7DI4NbiSxlcHVgpFh7ZDBDmWpxEVkd4qx
L5LXkxfXdFGmXePbEceShEeCiLBgNOABG0pKHcA2NKfClIDECBrF8A/UyOYA
ylUY+fyN2rzcAUgZTejNC/ikP1WEG7YIAidJH8KrRWORmKizPft0v+YfKsTE
pCmQ4SriEme+ySX9cJEL7sEV1YVtzwgfh7JrEaT3d0feexA2bIZe5/DQczPI
eoQIsgrAJmoQ4XvpoHo/oWhGPsFBePAKdVsmQPlRGPeEI7GGq8uWfxDI03ej
4sivhDzyoVcIWkr4CZhdElh6FEgNrZiKO1U4erY4+n7UVflomd4YHHy15huP
/pGcfhHmgweGAGSAl81sQHFiplc/v1GMjV5Z7vgbkx3yltVVMvvjGhF2rJvh
iStXur4ZSUB3lf0/Ck1nbJBxqWETbjbnHfVHeJgffNf8o6TzsGYTLeSePwMh
NeTyYAfwkG0mKKkCh5K8f4ptqdbP2llXwsgME/eV8hfL92P+diIhpnVgQ2Iz
bS4JDv0kmuEtMVdSFvOlYyhOqoIOAOKDsaVylrsKBHRjCphiCtw2qAe+jlFP
CB6nSQc5hgWA9gAyg1mgRC6mZmDo0NSMA0Obgv/utQsahZxnBRTH9SrU4xJy
mXeEq+3S1uu1TvX62+29wiLeBHu+S4C4N7vjv7mFspMmVhU4vtyo9njxilJe
DSYc00sWeovZ4LF9JEfb8vofva8tYYfOZRuR9Z1sUaL3xU0R/B4OlMr6e5P3
cRIi/ZIAy6g9taWRwZQp+7woV/j7OTwrJ1a9n7o8huAWfoWYD/a0p/8wwvQH
/qxY3Tg3rDjbTy+ydSovc4lU2DgkSNh9VHzz2mp2jVrnLL6fzul0X+XYxPB3
f94BDYToXO9v7tbKsAEprTte1tO1TwkL8wHGtOHn8ZsNoXDmvpM6iWUSBzLP
Gv8o64TzIvqebdlRuzd9DTKUZC2jqqcoQwhcxta16CB+DnrWI8z6s/AKa8Jp
PxP4HK1VrWFJdZnvtboZYsg1psbFLyZnkYht+9kh+2/ksmq1/FR0aS8glune
5D4DdVuS/cGuhW14uls2nAu7VCS4diDuq+ylf0pr4jcDFOWbLyxLeSsVzRpt
p+BP+f6Bl4GJpkbUiLlL3aVLHw5JcS+VeDwMIWGbj2OJS4qkb2jYUIrSi56m
G/lfQPwYkLtLLcOF/30nZ/ncwBd3rkdJDOPsqJzWM8PgX6lNL6qL2RDDLQ4b
TwYOLhuykfQYGW1EVnuA7VXQGEkt2I8GiiQwVagJwh3ugROY806Y+QEkivfU
jebk3eOaQpxDDI6Al79HZGgAeSVvTys+TFfSsgBpybKnkJm3AgGTClkgQKkK
KgPeL9cnrXHIOdOGWvfZmNUTHVyDEDxTydum/CZxN9ozHCbg5u0sZZY8O+Ji
j+8xsXg2WDyoFS7unSQSdEMHtrOz4EE7qc+Srb8GVi4bNowJFWr4sbCSrbDG
Jbsnzv5IptdH3hOXK7Cj6SBDWBlML/w3qqk+hi+WM5TSOGS9ffJ94jcuuXbJ
WjfZfffuUQMyk4lzPNxEHpS5KsqStcn7w5DZZjnkGZmbZ6cpHJCy714K5A3N
oE6y5ogfDU7xCw+SfmAsZKr4wVsnh0Uz8jbQ7TSkghCc4LeBWilcrp0eIKxu
OI3hSyukUrkk6dndBs3az7wyZ8shy7xyXAQ+cV6vnNXfEbV7x6SQloW8HYJX
oytZYXoi3gEHrhdVxlJZKC/3QIeRoVSXWy5KzO/bLcchRDfVJ3n81ksOaa1P
REDl7jfzLQ2mWXleAN0tsy3JrdnRvDK9/mlIBNWv6tcaFSemrkRal3wV2Cx2
DCfNJXIbWrEdIJIrZ9kxILVqhvLCY5oCrcKFhXkH9sU1V0Yd6rJzSdfT32ct
89K6EzuNQf1gYOWCeqjSYDXPvHxCW/96hoFlbvLNNjNlxI3aqsnDvbNUz3QV
byOm5EKDd5jMcQJR3oI+Kbf8cQboBrE5vwqJrmcOsVEnByLoEan6nn/fAjjK
P0h6py+T5pU4ZxE/kCUUxe5J1/Xw5J8kGBcvdp8NnoYuNB5Z+aJH1RRtnGd2
j7mPBWHhHfWFYYAAZsB2TrAWJYNysYC8k4P1tmP/IubjPy/RmfyLWGP5JSAv
f+s1ZXeLq2y51YmyljfwIO2nuwg63dvaYSdUG5ojSeW3UMPLF+TggWV2yTA2
G//Lv8QZUltonIkmZM18i8iyuGl6jkEQ9QNZneQPsMwkCs9jVP37HBQUffkg
BbeoWcnM/HDEt3qnB/rmBVSDiOZ2dFcF8XBUjYQdZVwGPLX+9fI5yJrocK/k
MyplFsXaG+ca91tyx94oaBkaLRgYsFeF2Enle5Kyvoewnh7dwdGCETiv3COB
LSlvUB1BjLUKoQnjOQBlME+SKMe1rOGBFpOadshUyvFs7hyxog70QSmzC/TV
yfnR0ap8OP8oy7TcwUOZaFwwuo5ju4/M3/LUnHDv1sHqKu/nt7mvGsxP1VPG
S11OQORTW71tlfw6I6tFUVrDe0KLhlCvAUUK4EBxyn72kH9Us331LpxJP59c
jy67mkSYrsKn1RhgoobdvAl35/CRCCWDbggrrZGgJC3iIssPVBiQR1nlsu2x
Hbv96N3PSH6HYhwFZEwbtn7SM9P2XUOleamAWTiBCam9AbydJLnM192M1OJJ
aKo6s0Lt6dFCPWeTkIprcREir/UiZYDt/CszNOTM3lqQos1VppcPxfvbvnt3
oD45K+zqkgYjSh1kvBZxBe6Cl1/LLxnlkGKa+4KjeChriZe4VP90pIG55ksp
JPuTAOnTFDbw8Mv+w02952rVweoAbTKGxpyTj+TQz7ui1QM1EAVttL2LRnH8
fwbUDkctc85im6U/I8rUncrB8hISlzKFDkmNTbfUgz8qShPjUP1APIROuotn
qYKGEfrbYlzqN05CntBt0Es1aPyMBmM8FqJ6nDqg/ATPbUU9wwFRILA28tVF
UDNb2/be3p0mazZvS7EWtBPKq5jjn0nncgbjPnk0L1GqoHs6W1Wzx5FyxyUe
fwkWCZy2QVFqP+hsBbRr2N8571rT09bsaBYfIr8hsYu6G1jstM6Bz7govInO
M/+Uv3dSfqrHiGtOtSplWFOZ5mUTLdZkbvaP1mlYjPf4ZWB8LVIBE+m6yeG9
Gt/LW5iTspKpyAS8Un3BTyI6uIdIn2eJKPd0fffmRkfF0/XO36Myh+pxr8/p
67SZSEd8Aq5iVLTPMUceH2ifCs/2hwnwY7x4vBN8jqjSkrH4eGIoAs7S3sur
g35QQIG4ZQEoA5Lxi/kJsdGS7RQUZoGGKEiRPPVOwpQD9o7XD8p5p8fVIYmi
EgvJFIDPP4FQHAA43+iPBvLkaLg0YMppEWLQCu8mRwxLbmOuZDFEpmVts+pd
FFsyPSDEX6NdDPj0yMr//vjkYl9X5U1bkK9+afwy7KpjvLXFOdIOWn6j+uoF
wUPS3IteO1D0a2kC9D2iPRtNasCE2lhRvNazu35rDjAECN4Ir9W7WNsJjFg4
J6rNkUycUn4zXGXmECTG/lRupr+e4zJ4ZFnTcygEkKjOujFLuABETiN2+6bI
ftFrL2ZYHxLNZmCc0VLym8CnBu1Bgdcw2Qt2tcNXYTGA5sQTXajDAG+pjOTD
D/h/7htkQMc15b9ycx9xLbu4F9ypJMFZnyvlBt23Fl42NRajhBOcxa+un6ic
cnGagwusX8yJ6mDAII9r83BnWhGq9T4u80ieaCkSRDkPoNfS/jXzudNTMkJ1
C+MFFROBBTkVWJe2XCmrDUqWh8dSK2GYSx+h21ktfp0pqiQYW8tzvln8SOx+
WMY8XXH0wwgZaYTHr96N8F3LgpCKshVPSksdZ66AUckXF2XuJa82CjW2QvDf
fFTbqafJcaGOxRQQ3MgzpuP0btregtht02VIc1N3Q2HWTipIHmt7AXkUjsOm
HZW69Hb8Jz1dg8IfF6pDucyLV0gYXOJcvQ36bZeY35HaTjTn4jv//AeNgars
Rp8jMHwfER9Yb0+eZ1EskZB4vYJKdbuXAx4me47+GaBoTFsCZtHOFdzhaGVW
cdajiyjVijUC5WnQDqrhGvZbqH4hIt+JekI6HXftT+2Ee+cuUjF3yqOD3S8p
pHcMqDH/Y6vwfhL0hbfSSAnINctetws+JRH/h47D2B26tI+JkwtcMUwLlAbn
kXdYTFEPFx3Ok+kF3z9Z72Q9UOP8pKU2s/oDOJctxikWzAwzKsBjPWvDu3Kr
ee0q460qbDxxV2F+/MH629Q7MgUrya0RaW8k98N/Nt48jFoUrT4ikQMWIydx
lg/b4ZUnIFGOtilLKxTevo46rCHWF4eZRlrH2GeNK+ufC0P+X+5iRSP1vzA7
0mze5N4e7VgYjkvxLO7ZskmFnK9MjAcYR0w/HS/0SjYG0faOFSWTp5m71tS2
MwkBojmXK5NekwLiLkgnzuDXALDJ6a2jWq63kyWkkw6q2vmfmvh2go3CRyc4
oP4dxEd5z/vFE3SocW9XYO1MJx+2VWw0y64iuM/QlubNLVg82osVv0xlkrJV
76laILyny6So3lXIe0uKcCDWXTSBPFeisn6igi17OLkYLCUMeyrOM6/adcGG
SINYyRhyOA3A/pV2j7RL8YRXcII5LqDglnRoVQ1jq4zKx4Y8+8Gui8jHOFPt
c3o4tVbp8jWHLoKYD2L9HVihJjuHeCQXbbByKL/Dd1SehwhWCNjsyr8gGUHW
wAdj/QtE2l1B6BzWoHj0DuBsoMq0twmtAqBnDcB66Xf0txe9I9Nf8tMNGSsE
hRTnr+v8HB+jx/EXEU+9MR9Z9MyszFk/bdzFxdXPSQ4anhurAxAD8oKlKvMo
0kxZCavC+uVDez78Q+LvSX8DsEdeFgVdFnZFEyGNOVaJsk4o05qqGK49SZuc
vI5GQx/3PZPSwz9MY+Y3JTK1C2W4P7grDPtJNRDiM3X9B7TJkRZK3MihN6Sp
3pyZg6Dwmm5V5f1HzIWjEZP/qWn69Zesb6Jybu26z4O3ZdWf/14sHWvNyIfH
glPAkrIt1VnBJESKUuEJgispkpOq9Jf23ywQwAXY1r3TenhKeZwYpW8p386w
jdmSqWjQtfmNXYVx5J9eC6RnkCmox9iv3JchNFyMwEOUzgMvIwhbuUgApX6X
dUSxTm/mkgCswcQr849QeRXSFe2Fr/uJJltwHdX+/1WEPfeOtbnJYGm7Bs7G
a+2zWLvui168QyZEpPPrrkJpKcpdiNgr9SzpLoBmJn9sYGaPj7y5ABQpGjL4
widuUDVMqpH8AoKFUIT15EQBT7B3auNJ5GVCH84f+J8k2tYI1BdYKxOUJb9V
4M8rW8VNXpmcsp4FGr15o+PcN5FghMjXoAa2wY5Sa+HsVJ+lvfrMlgPWN/Ju
7iRh0geANfIV8O44He3gtJLNCo5Q4fVjNKt6AS0wi+LOQo2UF1BOkhhvm5xp
C8qFGKJGgBrCAnchQ7D5wo948gpLgL2Bd29Ttz1opgEScZ9n1VejwlnlNts+
KlX/dJzGgtyLGJacmSkQ6LtufAEsijWXR7ICIek4tw8MoajTImV6M79OyzJR
jj4dfZwyA1sDWpFmGufrj3lGESAXE7vjtSP4e6lgd7zdU5aCyrQz6x98+z5H
ZzB64mbFqeFZFlceawRia5saybF0zm4f15FFC5NoWLby62LZ2NyfSy5j03Xy
x/I+05xuYUNZWM0R65sUS5eARFDgMbYynmcRKRMvslgmjOdEBfQN2Mf9DhCf
yULQUx2mBOHSGMfoxyar4ODr0FvRrHnZjPy/r+T47aVMAXeoDOWYrPXqtEDW
5rgglImuhzlrLpTDbTP8usr3qalM6+47K6jKwmWB7ffiFmdWwspz+KeQXmhG
u8dH1Edm6jVFenyhlb7M3t3INIDVIRu9YJp6eAzFlfaTCkLqdb/IbXG58jgg
RtMnDhvMaaxqBP+IFq33Z3dVe1L7vzeJqNojM7Ge3Q2D5/aNeEsqrxgw9bpD
ygFi+hh4sfUTDeo3+Ry6tqjdr4XqhojRz1zbcXWW8/mjMq8RmDmBJz33SAwF
Ou7X13tpUt3Eaz78lTqy88flZ11m0IpFFa4Wlt+EX7jWgS2JSlfpi/puCQbZ
o0xarIGU1ILgr8G0GG/qn7d+svyrNttcP5tOD6EwBGJZgXUAbA8X5dt9PzWz
guYX7EynmZW5VDtUJU13SmOt/pqcwF2qXZbEZeir4qnQjWkg8lY8qen+zYLC
Inz+R82jPvaZree4G1xHBOO1+RRy6Wjqhe9k/GCRB3Xyai3UM16gtc3hY71v
5xphELF2FH2NKNxxVAqrmDNCpqZnJYEZRtiCIDlpS9qMQrTkq5nuuybi4jJE
wUsP6oC/4Pf4MLe0cE6LqDvxsLmIr8GJUa1q+tt3sbKX/YX46nAvorfEhkQH
SW7nG5NkKBV34oBWb5EqhZwqzfSv/wJ7hAYNBclTk9zuQA+Bgw1H8b+AdyN6
uZKbVfG24UloD0+JHDIpDXxNWRVy5vAJ0NWs06bUoLmyHyyKr2rtiXk32XYH
iTwTYS6eyeAv+fBV31zWJrrkjB9hiR4BIgmoMv4yiymYBaxBkxaNX5452Sfu
88qz8YI9jj1Xy1igN6UiSMnf5ofeuGZw3qB+Kj+rCvkOmUbgMJnBnZqQqxZS
nNDmARoOy+C6n9y1dGX756snHPd7rkmL3cCCj+ciC5Pf4hjPKROVsGlp1VOJ
AIc6yJE+KjLpzWIXWSjyscIRs+ROjDYFiRx5K/ooVGD4q94eQaKMrGlnILq6
4BAgDrzJbXdxz7bg35LYQQZcAhNfsFSGLMMDiobL31xFdgbvyB+ynRgyuI+4
5dj0RoCdT1UAta6lF2d4vTO5TQizWke6l1T64Ll6+JOSy6ZrVoPKR4n8l+42
vHegGQFb1TUcfkIF6vkAe7hY1fcvoMbDAjr3GoFnSZF37IA+ubw7T2n/61la
XNYLmkDRws083SB8VmbBn+1++hqky8HLgtLHmbV9ZxIhSN0xg6x/IlfMYpSd
fQzaTlEGwwm37dwdOXl304/4BbjYMZqqlCKojtFBXuo4xXL3czKoP2GhYpVz
wjyy+Zf6dZxrHbJ8shXIvVRpVzhExWOAmPsXsNWDUoukUWCohd0C5Jjyiysv
JGxoo1hGixRjzMpoFyCWtcvgF9n4Ulkjh+NrPtGUS2vWwp9sls3UZBFCPELG
+lxdZxOiyEmYVyiQhrRxoBoKZLablQqo7KmKSXTfuvYEpJcMddiPFaasXIwB
FGEqYlB54GcpVSmxk1U7s8/303g5Wuz6SzuIpU16NpTtOXJ6YTGdGRwqbxS3
UzIQMcvXB7QUbUNopy7XqFJaZwF1g8fdW3OBgnLnsq0zANnbfOs54pRv9uIp
wsHSDEdpkgGccuaZhsvvXjrG9rzr9M1DdJ8AiaaJ/m9Kc6t+CflxrikVG+Oe
J3Dda1HxqzjiGA6DyaH7bCzIM2Dz2E8UCjQjRlkR0qVHgVAHbRvRHdyExWlz
9Bv/fue2PDlgmQ0919qlyBlqbUl+GuUHwcowFh9+jrRImemL0aWK6HdjiSGc
rq06S1Ldaed15tu1/FnhjmxJ32eYGAwGkGMb9aU7hU11DaQ7UF9H9Lw7vLzQ
LolPR8d0K9pwzQqNMqsxe1nAEjl1g9x++ODi2/YUUxVTqQpHwRiW/p/0Vykr
AUcHZEnA43EfLjf0ofF3thEGeCdL56zjC5u738EBe7vXMioAekdNg91VOl1M
gIghIBreahoJ/2khQcUVAXUOP6ytNE0U0yZ7xgLuPaLMP5OQ9abSVxj5AMhM
V9Fb85uQ3/ip+IBavHZ92bGx4MX0SOTt20rpHc6I6ixkHinMTmz/hc9NUzh3
RnNIIuvCIrvrVSW9pEcDHbMHkIEf2XGO+MyYEtYrSE42y2hqjzNMKEy5Xr/0
uVEN1akwqvORRQ8Sy3knlZ5QdJMWVEzw3MI2yWRy9nL7obHcRKSVef5UtI/3
PteKiXorv9G15J5j/9OI+9J2O7R+bA1gqxeuSM01ctIDPfcwdm7LkwMv1Ldt
DwbUYXylIoi+vSPykC6/MlZyXgxosL3oOuNuLrlUJ7TlLKoFBROcS/dUDDVd
M3ay+hxR4EjEkxMtaOp9HaoH+OZYkKS2Hsf3aBzgTp8xIEG8jWcH5WWPRado
ctMqrwOcG8ER0DVCqvvLLRmxNQ+0cb1GVm6WuLrC9qrKGlOyHgdHnXlfRzXs
FAYN35JXbmJjyi0ffmQY7m2+N0bY4zjo8spdio6nUbVt9SV3JpUwN/x9IfzH
xM06h2TYTMoF7o7qKnTGHbJzN8GHmFSrDNZS69vN+0+YIy/TjxLGsgT1iqcA
/TM/0sUqTDL+xiXdZ+Ce294RrMfhCZoSuLh39OiyY45JYujYnJSV+ymcPOBD
Cx143/Q5keccrGIx8sUXJCpQo92hf3kwx0NhELDJz62J6hWi/Usf3TrtlEbF
6GY0rniH1lBqL9u+Kgcssy8KxNvAOCBPLiMbRlHDJDsKWMBmtjRy9XpxJ4yh
iyDmuT5qBwsMCNLUpm7D4+n4GrC3OvsDCIMSCmLLVzPk/eJJR6ocbsRsJe25
GsCeX9B4zpebYphDBXuWSgB+Lz5MOtN7gtFA0i51vpW/QPjh/22vVNMViEVf
ykkxyI1Elfu+gQNY9I0MRcrUW68xX8YPoK6NaPODf+Jb7AYZTn/81Ry77G0N
xX5/XctrOLjNdGPBZqbnCgA1+deyMp1XpQWJMFfxst6+tP7WuAeYK5pIlBDR
MHo5Rqym/herzXim2+Pimza6zfMQuW7yrwdpbJ8PyFMHAZhYZEjfdd7gak3J
+OGpXhXJy8unAOKInzbp9fLRLBvQfLI2bcjVEyjHp9cch8J9hogL5+3p7y7+
FDqWOp/t5PSHxkuWE27Fgcxaw4HtHKUWaqZ/kgjATXzSFmGTMChkx/xAAb9l
Q7poYd5y16l1gyQJfqoWYPPRLG4Xo5yLQTjnLWJaUq1l4ICO7sUSD/bTyHVm
pkW7HTCpw5EuZZYldOT/exf+6i80F6rohXQRMuPMhoB8iPSHMmc8M0CeMY/F
KwGfuFaaKt3pTVWCAd+dOGUdVNX2zPCJQCsLBbZ10K9jvfF80VYuULzz5CUY
YDxQvgR0EsqvcBKeVCxqGFkVrfGyBPVL/UA6sgjUcY9yQy4/DPafQuxa33Kw
15W13zS/3ZTGn8GM/EFI4TSqJ/7MZebCe6D1fN80go3s96jg6Au+bqoYWefD
Pahmv5ISN4ZPuhhhID8x+lviN8cb4sevCaGwEIleLZJ6m9tV+nKODmw3+xEd
x7vTFWcr5vIVJs6RFKyzzCjVuhgK/u6fPIVm/qWhAIOyi98uore6qOTyNQ0T
c5MZ5Sn8HtshsG0hq/I/zyBPfZyCJ/T6uB6KqM9kGuTIhkAR5+Vi2P1kqSKr
gqnHZdc2ZMzdxLESzCm4ZbOY+1XCX5afwjjrAZSEVyyslNc/7Bip1Zemw+g7
vs4QjvyMBLmVbtyXKeTq9Cb+kH70UncazX4/dZw+W293uvoXmwk9JV96fO4h
MRZJyWrOqDM2Ddva7+KvNj5yDC3YurNIB0r/YvymTejKF9aYk7rHrKnYKM2l
I6UzopvFPpjIg5L9YTkOMp7H+QfR9AHnWcuH65dg3dvAsaRe594meIMMBm7P
4Fba+kdKJUijbh9aU+6/6xk0gGn+Pl3Qq4x8oh2Qqn3oOSBmhNyhJn9ZF1YZ
/Y6DnikZMdziS2JDx84T+1AoqdQp497T/qmaawG595HKG/JcPENfyKhvtg2O
2BU1CZUPDuqpi1CXba/wSsCjvyr9vyL83EypagTEzg7Lh92HjPivU9rTtqgg
w7TAdHyPP9tc32BSjra6/qhCW9WKOHymY/L1XREoZ/nHDxXir9upEmzxQQ0R
V2w8KCuUhSnm+jFTsc+b/IQMMPGR/RCSoosPRjqSZ+zi/DVyxCALVsdGk+Gh
aFj9ErMgqeIYPzP8fKT/C1xsYs3cck1ndcFdPgQb2R+g84Wh831OEgL2NzbS
T75pU+8D4TnV4HtOFIqnH+aPYITLCoO3JFHfxUH8ALOth0wpiMZwgIjKjFe6
F2vgENd8D1J76twGo6Q/zUu4jixEwSJkLIf5W04lScruo59jKg78ZXSDMiuf
E0F2euuMMSIBlf/ueccVKNCtDm4aIBa+ZxOjX4x67cd3v+2EFB32i82YxF2B
e2KmhAW76Bai1Oq6A+flmzMyLVL+x5vh4c/vxAAIc8OLirc21Qz2GYwzhGSj
DiaOv5WyfkUjKN74bNVn72Vc7tIUwhynViA+neHZB9ew5aF6iiepZMnqTdPn
c1Tw/rqIIdZmcjCskIshKLrKCINVLGcHQuUBDJllzDfW8w4DuWtjyuvTqzf5
H3m2R+qdZ9gzJcXh/p4aTva+kRs0UPQv86ONEIJP5yzY2wEP4Tm/iyVm3EuU
ChaYgZ08GSITbPqfmXQ9vJUgQGk9ydHOuDeSR/E1fUco02AA6rdUGWcgFSZC
VFjAEQP9XPjiMO1Q7i0RKqGmrPKR1uJmknbW26akHVea+HdQQsBiHZU36aTF
wQtlja4keQa3IsVyOipxymEZ5/bM8JPCX1iTEt+IavnqjJOwWOO0Yy/4iNu/
XORjDaJUeYJn4YU1j6S58Vb2pdmYoRWBnkRqO1SMhQ6hkHBBBlR/kr/SnBTx
WHvqmw4vrI3DyZkP8QIJRdMGDxtdyxF0Ock0cy/Qo5cTsV+ZsTODv/IN05+r
PTjhwqxk721/zcA6QS9CUhymWfmEa0MMub5GuYUmxQUkh7G+yBEKJ+m8EWvh
u/8wSuc4/ZFiq85J8JBRZwdM3zUGlkzgQYqgKVp709oa8o+TRrVw7AHMG8/Y
FhR0jbFsC7RlLFd7BQX6J4UYll0AlKuxLSSXEOldXvlm/dxbhosZtS1LMRYt
XnldMQZ4KejuQaV/vIwetrerga2tyWU05yBsKKpT54QMjRAZRNBjxJEn+jBr
3Y065zhapDXAz9RPFELAS4tSQeUzjR2mRHGMG8xUaXYIy0G1pou/QFN82keN
pkYxVAAdIVVvLroc0LHHevcOjJKeirbMmKGC2ND1ev3jjidjdboP6jnxrcGQ
vW9VQOOjaBjxl5rYXFLnu4uAXLcdkM322y43Qdh/sRnEi8i0toToCHteGINf
1UmLt3ayQHrKJ8bkjZJ1+E5Wshk5f6R/YQge3Aq2+IZIaXWADAcScLooLMoX
JfT/EcbCE00MSLQmEhSgO+KdDhH9Yd9yqdFaKQHxPCsiPhPAvqis4VGL1vNI
qz9OYPvUiAkj0Ty5QKoPCrzAXappJlfp3ll4oim29bUT8NBLA6Op7y3Oxc8s
ya8TGlNq3ZVXjIRcjQhu+z+rYOMvNsU+fl5R5lU92uvN4NEGvIJYBIoQ2PhX
yxGSNujNAF54BRRuxJNmAd9RxHCuu9yPJbPghPf4PqJa/PUVWmZ7Xwd79NBI
jEK1sA1iMZF22UG9mutBY6Q1deEe+/zncA9Vi2Bzs2xA+Z8lOhuJoNRDgJw1
nIg8MiuyntvP/yv1Ldrgox1/5vBCu5AYaWRgCQmlLNGnDFS1Z3GLeR26LeFf
0HcVymBOPaMVt2mREzGV6cpwXIh+Gl+D5mYvHK5esW13L05xEKaMuEJj8w34
G/28OnSsW9SOZfAEpazXl2CSbDpHivUFGpogsRH9Tg8/YJkzv0oxp9wv8rIf
Nvo05jf4WBdtgSLA/HaFUv+twlt8Fd02ZBjH1f1AHohNpMA0cmgq5xlDiUvB
Kwsv84UT+1+PMn44pPAUf1+du25v+wNKgw3pflmCNan5aedWW9cjFgGKGAUQ
Gd435XHcITiPLnarow+OsjTNCoyNvlmd6kmBdBrWZUB0gQBBF1vgAopNQ+p3
v3wvAlcrXDzh62FH1tayI4veJ98FdRdS4bWuw2uhEoRJRM30DkPBxAxtbZ/X
pusEypVSPlYgJZXmkJnT9RiT/Z9TSd4ApCO6BaOQARbbjbcwCw7XAIoN9xxc
ZqmozPbV/k0TyGISRy0nKJHl2gUMlPbAjXA4vY8Hy42pjvhlc2rQ9uNnd8rr
3s7GbMOP+I2Cni8aKqtVw6wPINaqaxKKpUlUisifg+WEkr7EAuW5vwuKlMv4
WRwEBjtXsG6oM8UNGaslq/ygdYY9utLqnqw0YIYVEgnqMpRQigqmj3V5eA5a
0VtNMe0/P1isv9l03Jvi1z1lEV3p4+t5ZarJDb0hEf0J9NAHIbTpCDE9yiIj
+5ujJ0cgmdHHllT4V+7y03tolfBPZQOA8TOm7YspSyiY/UnUWV6hThMr1Gxu
XijiPi+Y5ulRTPa64WirwV+Tsbx48QOJ7ARMZ+fvc0gXby/e+t85r2BNW6XT
s4556D09IdbnWhMke9+SjPAUSjqBZgFiO4SX35RgwDGoIMuuo7i1ugNXKmgO
+UB2nsQzn1Rvid6hZUnFZ/hLQFAbrf7x/Rhnax7jDJ1KawvV3NlLo1PvWm+B
1izLKb0nZTzze3SPDXV6SNrQA6TE11Ok54F+cMkbPxPVaIOyoCMeSvhjc9O4
8j7lcTizgHKtfyFr4q/oDghZ2m9MhwnrqHCGx+t6d4imTj/QaDC4cD8VRHGN
d8SdVJ8wWoXKwS+J/TdNnXWUjyMFEywwws8+PkUvdiTQW1dlUR16gY2VINJQ
ikZ5cYDTbJEv8QlZe3dS9BQpal9ekfwjB3TfjHgOaBZYN+GtvLOZNtavkLFB
LCkLdzU67FsIOmk8JmcDAFpMTWy2Xk4gF8Zx6joYgbqSJyi1AtYFbwfM50jh
0c/5Sdu/SVvYJm6Uz2rg1kr/4WhqVAhKzJ7ktipzIb+Kh/HyTaA9YNL+ojCb
Z03lwOHuKcQ1bpaOf0fSmwgGT+Ykz+KbcEaibHl94uTzl94TCtpwb/UwJLQM
eqCtpUJEb275+Yr/NYOL65pW+AiytndgZibcUx7THg56kHM3FPbvpSYiShVT
lbIttMdT/JZv5A+VxfVjm3iVPx0yqv5+Oft/yF+CVTfAAJOcA0YA+R0jznXP
o0CjzC7gkchPiWMCVodKuM1uYBxquPqPY8bj/HyNFU504nrhwhShmDfhTWOt
PTD4I3qKmO0GY2Zo7VdC4Ab2exXXdK7xK8tMTt4tuplJh/NMh3A3umFaz1aF
iEBSIT8YoUk4K5Dx4nt/qUPyODmAv8rNJNEnZX2ugI9p1g6xBmLIaJu0VhxT
OwNUs15EQWGJTdSAYcGojQWojp+Go/ScOmwOHsKcNTEDHb6YZx9hVkWoI/1F
afRQRusJmFRabJhwsKvQgPDbRjrCIVctmHw/IJT7Hgh5BRu33ROG3dzZ8Dzr
3hUqpgxpscoAnlbvwsL7DMnBWfB0P699V4LFgYKCsf04PybNyXkKHusqCI++
IsSSxPSIc6j+yfhYYWfH9j6sFyH7ifSjgpymf1Tzf5k08VJzyntjEH3HIxEK
XOJyf0KhDU3QKD8DfN+07a6vZXM7kgn0FK29JdIg5PDbXpBFgxDtoHT+dvtr
aqY/blgBCqEUBjuIljfYFK8z8bZpqXc3Qqd8zJrHhjCWju3PuSp1A4CyCalp
A5loDyuZ4DLIL3b5I5fTTqQwRgZrxV1t80VbuD4lAtmJVY5+kIqgIEoPBPuO
nrlxNwLBgxHa4TngwT0W71/gQhH+osxirP5PUqjGPqxrq2eghEnS7wNcFrJZ
nICG6mMMwbO3oeE89YlD13IGPi9RIyEV0XMV9jWpudnG3DDO/eXr+nD2McPh
9ZPzZiTtriEgvPdfPmNmP/0thbWjXMj4p2etHgYGaXUXAwj2bG5DIHHCjFT/
fX5wWhXxwjViUPF4fmj5v67gT5qf91Vk40KgAbrYPy4o4rCa995uaImJ3eO6
vj3sk1ZtyJYzwke0EOO2IbEZQEP+EB6b6gQO2xyEDdbF3tG8R0aY/AVwHiic
wiygjhnvo1mPeGIgiIJEFryQFUvLEeUeFYKjLZBZ9hyR7huePct8evX4YDNj
E3Kquw2JJ6QVbKCu49DxzC5k9rWn2PNuv1ipTBYQ9q9PJbhYpBJaJU2d2Vn5
3JlV/n017NJS+dtmZOsiRZw0dcoxu9ep8bE2tVfy1PsEPlMffWRyXzLb+9GG
YnvZF+xKuAbsoIqGVc0AZ68fB2ytSAZUfjl/6d9QHKdLrQKtV3CNpXs0Kex8
rDZTASgG55ZoOgEtL+qwZA9dHZzlYs1bLq2qYAHa/BZyDNO9yG7YUTvLjPe7
5DcxsozuFyt0wx06e4hiGvLfEV7PIttxNXe3/b420zQ1ChbqfObQMqzfc3On
Tzxh7OnRL1JpChwetsD5dhFwPRq5IWTZ7dnVzIGtmoa7YB7Jg5syclknKxd3
ECCGzlNWLW6d0yrODJTjX8OkbcSS5Wkzq3CWihmjAJTYiWPk0Kdeq8For1Ny
xIdvS6KBOXkxTo+mdGVs94YqZ36kVBqDUsidOfMF4ldofdA29JyimVl62sFi
5WsN45LSvkQJTuNDbHeUT+VPQRMH1DBEQTfc+nG91KREeCtaTkjOLJg/ynNF
O/GRkLPz4e1wBYCJMSl3QfzO8kr1ykFBmmi0wp+2/rHz0j1H7G3gFHAlHpdW
7aLszmtr0a+ocexYWDlEtpynJGlMsVZ4E0xp0Hg/DFiNnXQ99Uc9ycjqsjVL
IZZ5zSZRBriUql23oGtbl7jHha0pj30iq8/0CciNjaS1cbSelc4fiPFYhbPv
p9b6mShrZCDUJK4mx31q92xMwjytRcJIKe0ToAHeB39/HgkJL4XIF893Lf0S
y61Q9m5RLC5KztSwVRqUdXIr98G7C25pXkhQVDpSMDRX999nW/YBLr1/hcr1
+cbXfhsV00lgqfbG/6aJ6nzkZY8cS61E/QvfD/wY8iI9lrpL6kzPBXs2n0kG
Xe/7VWOS+eQwU0ukL4hPdDP2dyDkBPz/8qyFacnczLPFNr1sB+KjWMSeg618
c1hLHJd9CqWo7jWimLSYk5RPMt87sWxLs3SOzt9NFsujMp1dYMm3O14kpvnN
uqlkXq1w33Ht7/xql5y8uVuyl/H6Xv0zxkBPyFo6okDrpbQo9NlOEWCbGuGN
M6DYsMNx+9BqZ1AQT2ljsTgosZ97sX9a0bATj2IseQwqnZIHaoK1y5bnjITh
/xF7NuNS2sMTdF7oqadtNk1hkfYScUpjjagdGroqBZLGS6KNNSv5ATb8Ka+e
jGDo7gjXomGKfX+OdE1m8UpdhWt698v5D/pPS3lDqp/dZK/ZTOL0qEl1dQhD
NPFVmbMVAjkf3eQXucb7N051IxFOJm59I+ek70uDLnI8EZXPDplIEYDcE8Rh
+PNLpw1z3xlZE1GWCMMsZ5HL13uqy5cwmewPcGWwXW7KBtFY98R7zruYeMed
itNsS5WZnjXFytnnzMXgo3V0P619pcJjAWK3cwogBxoUqK00s/U0CBUjGJn4
aELIo6di5soyETyeRUfTJ9O/bQP15GM9JLz4ThmDCbhLQm5v7t0UKCDwMiaV
m3rz5AdqlNsouWZ6dfm+KZn43pT1b9J2abf/Dr+r+4u67ZAeO4OhSTM22FNC
Ma9Jv69D65M217QyXls9jN60XCGP53P8T4v83508db2nl0Qb6g22sIpwJ9/l
MxJHHOmt5+LTsC/CD0Afr+YInJoNlxaAGwkZiYcZdIMwlUqFD68lRGkWeqzW
u9WD+n3UmWI6Lg63le/DTHxom9cxhvKkg3UUDb0V0KbZdGJTtRobwsgkn6Vv
WQKw7WiQQfpu8ozjXQ81mTGQs/ojxNVMToBZUL+gF4fhktkubLP/6gDKu3FX
XDommftufo7tY4Cl3fxbgWEcTNqMorWWXGTxCJYnnyWnPWiPUQACnWrnQPH+
WA4JL4bF9dO6dXUQSJbTirhdqkmGtvqRPSrmVfPSv2MdN3mb6tpWxD6AE2eZ
6ggKM9/auu3mEOoFxX0mkkOmKSGzxxNYVqVt2HvN2CG/TMZSjiCGAUmYa/jL
ZWiIniUEvIE0OUENreoyv5AisV6JsduCS4f+yTRnITMku+Fji8gOi9j9hfny
VgjIhnb8/LIYroSYvH79575u2+w+b+Afj2PK6fHmcZQaG5yiXn+GTcTgnQXa
C2jS8J3PRajZwHe122UiFuPkbd9zYvJ4Sfe/BQY38iqSyee5/79elInXZ1Y5
CnQOmcP9kbp7wjnpAqr0ff5La2fWMs/N0xBp9SFQejuZEAzrSsuvcv6BUt/d
G2A7bHH5kxMHmJ6/DKdCq2+T9TDPDiZ14mOGE3Gu0HUb9VXqCZDRiUZYB0b9
KfJzCX/eL7BVc9EuTkHwuJAnKWWZGKQfBNSUe0UtqE/1vOk1nTUxk47Y+7px
TglHtoJdkFBoiAJto+zn+vyGmACtT2z94CWZK4cphmLASivbz4/3lwACKtPY
du/YoX2PheNuGJJDMofsiUsR/XygAobOkljuljPLrNCroFcFlUkbqSFNkGhw
izKkv34pimUYFX0QBit9kWsyA7Ssp+hkh6ufHryS2WMvoPvke4slQ1/DjkE4
Y7gJFqpuMwinJs2//YYEWHbNUKfrKxLVmo6L3/gkR9oWwRAjODewt/E7+SS6
JcxHEGhUKLNnM4TS54jgzmFx0Dne/Ei7Lsyf6l/rs3KHaB6KzU7LhkIKMQgI
QHCZtIl/4kW4ts1uj/6sjomsclxk63ZMciVEVmZ6Ut2tiTlLtu8GlMNzhj14
RW7rKWzaekvCx9/A0MVrrNakGH9B7dfzRyli/De0+WYY2WZW4FnM3hfMVRfT
En/dT8foodlqnDW3So7bFkLakfgyh7x7IZ7GAZWVhiwEWIKY3TVnwNPSSjfK
IJKwLSOrwlPL+jDY9BQtevBRx88JeIR7CaJrLn0qxY21p/DyWt359+W1PpzO
y/5bc3vCj8a5ye5BbemRiD/OqvG2PEMjMCsgw5NO1CvW20hn/wJ8rD9bS98c
gcUSoqwajhpVZ79qvIdzWqmqWb8wF+3beMnG/UVYakGtaPzZKcmrqP/pqmN0
r7QObtVZCxmq7e8P3exa7JBvjIjhggeUlfv7bUhiIgKWi2m1uOcRbxqRqngf
NPvcttvulQH2FGAp56hEhRXZvzeH2MC9gWhCSOwIpIuK+TNLI/UExP8I80CX
mQ9bVIH8JRr2IBcGXino2pKsFLSLJ/dWTWG95F/yYOhmWl14ralQFpnJJLR7
+aHcSudOzjtrh2aaRpifYrU+qw+i6R2FHoVXQzJ62NH5/WTjBB9nfjI3r7tL
8KyNIcPDM1kb/oPJEdfjQKuvqgJPOMsmmgMsKc/1cO+E6MPj/vmLgoJSDjyW
rxP0yLyUdubZt6QrVkyuNUD8560utww867YRwCkbkWXm/6H1R5L+wyhhTlW5
VZ2ZqkmgYjEBT/GVzj7kglPOJDmKJ97yQjfazVeDTpkXKWDPWTk8Jc3z5QsJ
MRpf1TMjppQL47OrFNFh2D7rp5ssDlweVUOPm6W50ysA7VWtp7SmXqMOKhMQ
y52ThiPSQ9swb+UmKWJgQQ5nbcyiB2gVl1XYdibsVwp7TrZ+n+a9Ysie75Nv
WPf3LiqPxfCjTB8S54nRriYyVG1VlgZFFBXHquammBn5kBfWitN3xXDHfsoi
Aod0AZt4RCg+5zRe2X2qIDjC06V6Hg+xnhHqkGZjBDjgG7EZ++HXEL9gXRUO
unsSWPUCacjRAX081NB5sYgBPXN4rr1LJNu01qMKB+k8zhG1JkVnEnnUKz2q
uM060Y5zFmNNnaNGtXmCuRLM2HCohndJaQtPG8AwsBs7VEnULiAlRsOO768G
avrwATspiSmTHszOpyscwgSJYsq6qd/2bbnm7TMq2sOy5KhiJ9GDlty/xGxF
7ltvf1qwJF7TwLcIWb+ZfDyFxohr5xCCmYjV6DUTDte1SM3sQe8wBucd+LdW
moY9YLkxZOzQfflzsBFEq0+0ptoF4YdtElS++fY3cM6h0mjfmwdcBXPDUOVl
CoYF196rlEZ2q8WFFkIQP2TrXAwvXRONHArxg89G2pDUOXLQi56wP5whPE2T
QiAIzORQRBAL1nBo5N6T6gDZQM8uJmrnNyFlc3PEH1wkiNQvdW4CVh6+PmfH
4gWM9n+IbqofncrrTaOP/dFfT8dmouE0V2n0nsZrkN0Ae3rfBh73SlfcmV4N
DQeDxkedYoV6Pn9OmCxsOTBf64ISJLRno+pT0bXs1Sj6Ho7vWKsnGTEhCdNU
vvjIdhouu+Aw/xg6Ul+h8/ArDzoS9PPAguS5BtUXdAPTab0oZqY27ne4vznc
ZnyVoB07a82gGk6Ci2ZsxQRguIvCMMBW/9USJ95+c9bSVMfFzWH63AAK/DTe
1hfVv37arUJe61ImHf77dHvOo3QAKm3Gz8v55XS2SIcY0MJ1Ay6mFklNKCFb
qoBzuKOv27Tbr6ARuZ09ubDNqx9hLUMshLoLxYj/Wp8p20XAByJIVLasBCCO
ttvpfPtfC9Qw/0qBMZV/Uc+6j45PWHFUm8PH+7+fIwv/zBkOih30iWROOTSU
yd3787/1ymk0/lFgPrJC5ZXgzML+S52K1vlgG9Z5iJ3Gp2HYAPm/LXnOAFfx
HcDt8O+/jdyXGTKhgYavF4W1aHYpARA+smjeWfidcO69erM+mLYDDb1vTmo/
e508hFVP8qUduKOzJPM+ui6xlvMXiEB6xuPg50H3515yhj+B+EpHDPlw1pf7
tc3VO2gT0V0SiKdzIKykRbFrqVaoTnpC8dDknaukSkrlLxFvl5PMITEw3X1M
NLe2aqnPVGeysD0YKcgjifuPWvY4GW/zZ7D9dgHFElwcZq25smFEy/TlqyXZ
ZKjHEsA1aHw0zl3vbEENthpIRFQP3lYVCNQS814EAk7aeqQg6+VwtXs1m/+v
PKzQKDNTpYneSjs5LaS6hlO3p7BMvtvziN00UhfjRf9fSzn7V4yGEpRGDJhG
SrnsEa61NQ9u/GOluZ/vDtu7p6tT8eq3Z4/mSKDjzXrhPC45mQCe7z+7vsxg
rrxUlnYvcHSpm7kXK60sN+v1hS+hbBgVN6GWIaoKcPhTNlaaIzWupAGEjkHk
T1O7b5RYkrsfbStL6R3jezjVgAqg4Xjdh+88B52Am7bBa4O8E7XJaiBBMed9
bktV46wBc/7rbvJyOf5XW6SWH0Px81CDocLJz+D0mFzcDuuXmMW5dVUnYq4d
WuF0jqsSRBs500Wiwc7CnF11zBeKAS/hTnyoEqmNaGi9Ii1fHEY6qoZhpQeA
1BbT1W82iefOQZJq4oQALMpHeJVmk4oH2Sdde+JeAPJFMf2xNyL9RJPwNzm1
95SwW+YCWt3kqpsmc1lfdg8fWeh929zjf+JjvcODnCiu2ve9584n527WoYF+
dNNnspmEXicA60Ms8I+jOTjMnip6RCXnYrgnUoivXy90OY9p3q/q3rhGp8vR
L5HwIzCOtq+rZRPfpw9hn+C5MyXZ0jjKjxIUQ2n9Wp0Bi2Y8V/f165YIrzqO
+344P10A+gX0uuyE+1S43m2iWTWjTZoA4znurR8uNWLq0/xBkle//LWMEJrB
TwwpVW01R7Kh025DcaZ/LSFWPM5m6LQzognuOuWQflRybXzCXyxbxkt8K84S
iTRKLdy1jvKXBYSiwU7js3ZtcwyERe94sfbtPCH3HJdwFlSVG8xCWHLY0l3p
9reFZG+gHuEXQuE7Cy+b7fXNVZaucGFIftbbyIx3S40z473vHLua6u/v1oTc
RwBWg14wg6yWfp18ZjBrT6RIWt0UF7cW5Ta1QdVSWtmfJB2nL6ffgIq+kV8Q
6ZipvoEV8KdK6RxIyNFMaxzCJ4DK2It2QQkegGl/vf2ZaUSS/c6QX7GdtFHY
X4w3ozrcrcsmdj0YFvrrO++l9D6DpKi1d97JkKgJuA1Xb7Imglzrh0Zf0OEw
OdDYphEmg0UEg2w8CMtZMCU8SRxuLs5MsBBJlHF+oklbfFDJ+INt6iS1NPnc
tSYTYkx+ewQbM6ok2tmcm61s4FbPbQq2C/sDIfCWgmQyCaJOHjnX9srwzXw2
pK2kG266NzYOTzsgXCnEecKIjjrQvyfyWsqCyhwRCF9i5L4v3btPAT45Go71
3FSJ/kP71vac07s/xkrVIpMEDHod8X+Aj+Dw/Il1wuITHBNWkJxQCa/3sTpq
vcfsBkEio3srxpG7YPyijgFGeHHkibrSf45P+5zBPwJSNJK3uYNknsGuZBLX
oQa0W12Re3WF5cPAjFEwmJ/SAscKGzv9hQfIDe5QMEadkM52f3gxp71mm+zP
apWVtzHfs0QT66dpjYnxZxsW9F4TURZgDNmTKSKR5b3fmNwsWSK5Rc0behpl
/ettE6LIN6o0LpraeNTZJ8MowJpWDs9TzJm3Ub93RdPzB90Q21+0jasubrpw
U1jdaz+E/Q+15tqIAtWmQhue0jbDnUEk2rHZWxajQ4tRrKdsl442HrwIadmL
8U52oI0n2vuZETGAwwUY2JVsi+lc2anZc/kpn1Q5Msy/3n1sx8N5vHl4GlrT
l6pOsbCxI96LeA3xc4b4oB3zYc5zN5hzR93FXRHbd9m4Olmoj+847xadZw8/
LFNeEDSvNRGbl3BMkjnoTilNfVlXptbx7BL2RPD/j3ox7tEjEPPLREBJvxSj
nBtuIsQDaBZcXrTLzVUdfh339WyPW7r4FLtQ+4NrvunMKpo75EYN+dvo0/hD
kiIi9411j3IIy0IfezJ2oke5evsbVPvOzsAWkjeavMne72ApbQO9Jz6CcPnt
Nzc4it4NPngnLNxzxAr/I8soNvYZnGMiLRunJH+lQkQgM7SQs8fequFrCNOS
UzfuyjChWESUnFY6ML+YSo/D8+KQijlGEOps0gSyOwmKKY3ReT8DyUHo3jMy
O4/Ix5RoXuPKSk/g50Qp5e3QicAedCPuN5KNkgSUdR10nAtARXLCBYfhpYqj
Z2bx1f3wdSDu7SFHxVy5wjsU6hJ7dANIVj2hTEKTu0BQMZv3S5ndyKWMMXAm
WLUHA21jCjnH4r5BTT8TBJgKTNh1iCVldKkVpOv9HmwrPn8mon0JQDnGKIQX
1P+S/UVk+ipBYWRG83vIQLlgv/bY/PnzPYev9m50VCyLISu2AiB+UDeRgru0
Ls4nfJBj6nVmINU2LgVk1ZNO55yRxP/AWRMoFfTWe6kLZTTN3fCpDLkpf5s0
DHUFySYhiMJF/sjx2SF5POJky1o15oY8GG5urtgkcAOUzbPRMYexxHFkjYqp
XR5b7y/UmjC7MJvbsu+tIZ5scwIPGLfO5s+IczSxWBFWwM6LGNfSEL1Z5ze5
gsgaeVhcyN40rBD6WCuyZw533wEiUZx5yiJdxUbsNaRIUScZLD5cuhQYhc+Y
LmCVJycz7rEpwc53Yj6uX7XtyMGHZKGRAKlKa7hoAa45lVj2PaAVa+p/aajx
nOWuJjWl8UEdAszWaZSvwdyrIxbUPWOBvsK4C4dwoRt1sZQ92J2iEX1W3c9k
LMnWwXUsT3uuktFKJNeKvJOQ9S6DuhbmE7UHe+Bx+mrb/A9NYk2xM1eiQsTi
3ErbVmfadOXC+UNrZ3DeOkSTldJkLpVALP+x8OGNS91Pu50dAEC+Lkb7sYNz
WjIdSw/WUdWsAYZPPU9K+XznDUV8WGGcoPeQHlw1mJXXW7Qxws7WkfDYdxLH
2cdXxKbEopojDI6LoJKTgbcGBUZufwdLlJLYF+rAwgx+LCDIIoPeN7lNoYav
g1QiBAgw9h+yZurr/KaREcuqQiJ6amTWnsAle63eKQMuNgeVK4mFAhpto0IC
oB5DdoqexvQlfbchIDPO9Yf7Fv4FXUXJg1rTvH2ZXE64hqUL8/VouxB/9DVs
lo6CrYvTxPlZ2lxQb1uqO4hQB48czTtkgeyC14kMSDV9XfMXGqOBC4WdxjCP
+ELT8YbtIaF39sLpSpY8XJkOef40Hgjr8JlF1xsOzXTq1OGHRwqasr7Mzb+M
dB6bdJiNr9OGGqOE97/GERhF957FJUvCCbqVhYIM6cDmInEFbMY8Lj2pkaFe
T4S2TjsDxhxVJl3tjRS1H+3/+L+0pyBNOu+HonS1OYbXFzw/uIHRIcqnWGds
z0wGVjiBTukLC8obzgzWoJJEhH2iW2QBLA/G6Eo4rWba6UgGWunwXWbkyLbc
Z+hk4naLrc7eb9OTkYvmwrhd/u/DXA2VTeYoY329FFSmOGtFdwFkligyYLlU
DWbOLYlCX3TthptCuBv3m3hCX6GiFrrXA2sa0qvz5ZuEbEktfeOhe3qSrndb
j7mI0UPK1CxGNuglzoth4k7pvyFUkvvzLBf1TzjPdnAkUDbxvo86bP8Rp1/T
jx9aAN4j17KHKse6I/iaobxW6BI8PHgOH/zn6OpDaCEe4Kk8lxEOvDGMyTkK
LjA63878hDY6Dg2b5HqIsswIRbLlPowoIaG/TAQIW0iz5S1d/DIhyE6pf1Y4
uMVJB0mE8jx8PaJBOu+3Y0Gxdpq7M6GZEfyHh9N16/pUGKvscmRECgkxWNno
zGdIHh5XrzVMaTdwiSei7xkh+osPiPX8bq4a/C7UjA6iN1lHcr35tlLTD/Dz
0lwKcQPe1qKzcETeV4wcoMbqqDzLAvRhw5npkN1cDv1Q2johoU38f4KfO2sE
TVJcDZnhM2lDEUUnlGrpqq5Q7X9323FN5XrqBGadi4odl/Fpltxf8KkCsGgC
SZ0V7qDsUqvQ5wPPAc9qjLHikHIrAi6jpKY/wUailLywHYWTRxy9RJ5CiB6k
uHMlNo/HGg6fzTIKGi51sAKHPufZHcsSm7W2UqF49iTKFEWKrLY+mFC27Sbm
L6WzGBaQlaUAwW9lL43eTFYjZg2QSiwaLn3OWigL1mx9dzmU5jj/AXQCGXKO
GEOi8S6KG0rk1lwglQwc9AO3nSD9NfqcAocYv363v+dGr8Dx4pBMpU4RTVRl
ReHdXGu3rQUri//RWfFGL3XsQCUPq6KsHwWdUmb8Bj42fmqiQEtAUjmaA59Y
OLFicduW6JrI/Sdwkan0V67jxfdGNMOUAMy8R0zmb2+cMQHyHhhDR8dLLp9f
HHu1RVsD33SjxI67T28yUW86OFtWMdFA9wIaeHURsOffQmk5N3j/yty4hXYa
l28KTHq2T+JqBDbRqB0MAO6TQEiCfXWpW722LUaebvzc6b+Sce63dJLkVwPz
yNpPWb42RivJmkQmddAjiv3/lQF+k9IdEnkerheFjZ1x9HJL9Cm/28iHi7sQ
jtuhqNPSKpHwVtd7UOrQtQw3nYkpfPHYBnz4XtiF6Rgc+P57yps0NJ8kysba
emz/AXbwb7Uv1X9F3eoUcVN+uWCJahq6q3pbBNnmfu32SA+PqXBFby1LkXbf
16rjrea4ugyJh5KNExakwe+SzddWUKPh1jLQ0k8kXJp2jTkONAhCBKRJaAv+
iv34y1SAS3N1Y8ez8pLa/XEaziDqOJsfmtvdC19LeafrWqV2ygc0lk3ywKWo
YeXuZOQf9i8SIH0MvGXr8Y85aREoC53DSYC0EqCXKtugm5H+1VaLOGE/KmdE
mdalJyzwDmhfa/tqQVLkAa/ez0oFYGn89QgkUXtER48ecaDa9I8FJJWaHc/q
WIbVFOXxmSgu0ryuwc+zE2km7x2g7D30p6277jzY9U4Pc0CZe/fzfGPfKI2D
2crOSzc9TAuwk7pBAyWLr6IxiPXsBcug//vkM3vzhU7ruN5KvamVpgSoJwUP
9pmGScFSdwBGIy/xgqrmvEO4qK+1vxwExtsOmsNAscA42vXhu+VrgASy2VEK
MIK2WYu33a6eKpLevxzBlXPFFhOIJeb/VKgmGtcDmsp5tHi7IAjb200RM7jb
y4tNK+aCaLcZqek7TeHxBYIHuW7cKyaHRRxoOqGmwGcitYG3qu+P9xhqodjO
daXfQn5R6zCbi16lKprXFE4XLKNGJexGr0xWWzjlozEqg0KLjXs6w5FAgcN2
gTaq5iszVtSsuZJKB6G34xaZcvChqwGMFM5hX/ojr3dXj31S8jdWB6J04Bl7
zFKYYY22j/AcyqB6YzfDta2fgG/x3J7Qkqr78rQzV7LlKjkY8DNZzJorOLfk
MR3KQEvnxixhm7Kil0T+OJbV2fw8eCZRAmrpZ6DCGYs9mbYAn0BrF2Rp+jI2
v+uZlJF0IwIQCbyXB5e8VvOcxPpJwHVUeuvRecidm/QDtPbN+SrC3UkelqSP
1B4DPzVskccPmTu+DAfS64cOPFoFLEiZrzDHbyYwGbEuG48H4C0IyWZ/q+Dd
nKYo3SDfeN9SJziUGEjftcZrQ+WKd9aj1z9lMMEahub/kkk/SqykivoBEOOY
/H1yPbr9xF2BkDvN5VFscsbZAX4x7/E4tjIJHgcMEObNl4BMyi4lFZYZe0XJ
TLguyRCjGbF4zPwqzw6Te1BJn21sZgURxlTC62IlPWIP4QYB0AlZR1XnQ1k1
LvP5xtAm7ZwNMWw5LrLhg7X9/sMSBabprUHJtiDp1S77K8dLdGfzV79r0+P/
84F/DePHUnKaBtQxNh2Z5MzSxXFLIKYKaI7JPXogM+dMpkuPKPBhN2IFYdkg
9P7VtNCO0kVy+GI+ldRdlYKmNinvU4hO5SvbO2A8UJVR7gxSiYOiek2O5jdz
B0WQGZc2sJweGUgA4GWY0PgWkjZuwwmOI2t0eZMaB4khCdeCacduHDmPIIDp
fPvC7+QblznI7+atSAN7ZtZNlvirvp7xgewJB+21TEYCbBbruIo0mRGEO+HF
5rOXrc2FyTN+TmoW8f60eVuomcMAkNWkg0XiP+CY7Fb9CCEMM23FPQl+cps0
DfS/ywYtplGotzm7qtUEd4BZL4hC1FMOeP3FgKNpEaaZ85MJGTiQ6JOcHJNh
+it92oCjuQguqo/gPL+/If6wbm++UMRAAKdHDG/0Ojj0Pv040LikPtprnMXl
ORYitjtVXMoanf2T0Gf1lip/kCfU4yFTCAsgJjdI9g4p0SpkA5222QdyL4RA
di4RX7TCELG3blkhr88KPTaEyqfFguANnOSaUFYXBOcQca1kegPUORMiXsb5
cdFBDFNY+pahicpzEZR7oSpDuYpIcKpOVprvesm2YGzDPENqdJqUAkee0nHm
6ISh6k8jbyhUraEk2dBd6Dbt/XeEwkl/KrXU8YU2GJT4a1PDGVV7zxXVXPKy
XfNEXwX99vVHFbwKocqbsBHwLC0MSF6JVZy62sjCw78nmuWG/iqqivvM1JuT
a5V/rejnGLp745FnHWo0U2w/vNiBcKwwQx/z6TmNS0sjHdO3V4L7gJ/vxHXC
BZ8coMA0NAHg7h2RwsPVCCLf/f+l2izcCvKcGxoJ02Imac1OzGYnEVyplPqh
Mq3tgjKXElKeqwE0ZjRdPs0w7TYzkGuYoTdS4K1BrdRCQiKHXIQ4xnQ4bTc8
JzQEpa4RghNky75ymIOrS29epcUbquVQbKMWmLZDyzh6zr8hjXx75SqFHRYv
srehgQT0jU1NGh2FL/BMI8BCOnOfDrIWWOSIQl9dzHN04fdS49Ag+RBlVzTy
BR/wA5/rO1xvviwek+7Ot0DX2of/1XrlqsD3+jPUGM3yIanw2D6zx+62Bm3F
t7VKtYjUEwBXCwvONFIFPy0CyEXNVERY6lRmxCOBzmF1JyW5Ogh1ZZfWD3YI
FkVlDhyS+BJm/d2MclbMQo6VUQaGwscuGDIAsVePWDABYm9Aek1SQy3tQ5E0
j/oZofWEymoOG0mHdpAE5bBkeqDciPtF7eptNGCUGnqynKSGZfHgpPiv5LQb
0o4AfqhROH4EKjg32YPGVsll9YzzUDyORFaB5vlKYpM/XesWGdbCoggTJuG/
1JXCPuR/Sd6LgAXHTACBBnJKdRnUbl4T+9nM4L49T5jqRpB5/SNZz5D3gk52
PTbykHqD1ZJTbS7c60HRSzbnRGSwmCMCKAAlLagtgUoSnLuyVcFyVi1doY82
sgfxWdykWzovg0P1DcKrUnhQQBIOqOMZ4rc7x3F4xSWv61mbVw9EZHPFHKsy
2TmP07aG82oYiv2p7HbpECvXIaFnBiJG+pMmw5+qGPCCRzy7EeCtTkzTUxOF
80u/dtOuqWDMqQRM2q9IZMDgP+bYI+W7l+laPaKXwsP95hGIxUOJ0pCNqjrT
4EbmiiusztwNoOoc8ziYrV/cI7Y4MzG4kCNOCojgow3+zzsMuchd4hu0oNg1
i2fPMEGh6DRucgF+iVPOXFC9aMPC3Y6MidGRVXrs1YYIJf3fZx46/FLNMfic
kkRZAJRS2LWenLXzsekTDU7N9dPwrJjaol3znBX3//Swr7fW681iL2pAJOPB
SEjDPyLEC3A66gWWYynPjV8p2ZMkAasnZUdjYMaTrSxCgledcCvva9rIxdzJ
egSTaqJ//nN5VKPC+J76HkYtiWGLDlInL74mad9ouUdz8FvpsQ7UDADnHplt
0ch7QGVe8KkSzkI9AcJsXBnRgupFDtLS07qta4df+fG7H+yTUQZttcPukp6W
K0jhQAA3grYSq9nNfI5uAfYOv+/hsRvDVIk5DSRsCX1aVVptA5WOHDqQofZX
pm0GjRbO+z2xijyjOr3EticQq6+MenHsF+IsI6vH+4Afhmx9YW+Mgz+Ff46t
juGRENld1TgJJAAw6/w+m35i8EbvShzVG69KMfw02zetkVH/iS83LoLhfhLe
DKRPxF96VXeOjNc1C//Jc6c9q6EcOQwjZnedxmYMbzvaziGR47NVC3UaopnS
AHT8WMMdFdgw+Sga3LkSz9ooJxtI8pmaBYkY2J2aFWp/tsXoKJ9sgGabBKf4
y1Lijh1zQOc/O4IeAr0IOt08SmAt2NgmJXEGZfy5uubwdjQJZ4rec2HKThO0
TZUTPrde508/m8eU9TtwNrO9VjXT70LvKHQzp2TlPC2K03sOY5MNRA7IIPEO
8QjK9SgWUCU/iOJjj8IdaqOp9KlHeKZ/AjYK5E9wi13fgIArO9BvfRy7Qocs
6R2sGUd2TpOhUIeAUnhILlfX4NxX91UQsJy/zw5/JvBuiyCno2vKyJDOlN8+
N6+K+yrO33/jeWko4Y+m0HA3wYOhqkZTF4bqCs13yOP294RiS98n3aiiyT5z
vaRzpQjwy8wCYDZTih/10sCZVsNV8z7QXIytdKENIFdV2OALvY9ZzhsJWb4i
onfiumT3zt0aNIcJq5SiHUfPeta8TJyIsajdx5V8L7GdiUY1RXmg7sUJKVBr
2qrwnKlbp8txIdrZoH8ZemijY5oMZA7Rfapqg60bY5Ha7MHSiK74EG51TTuY
8oP8Ky6pFj0/5mzaeZjBQJKt3mqORklpd9w9rs/yc88ZTrozkLVEoGO5h7g+
aOyVsP1HkpxsvbReaWUMpb9TScZzWnGOBGVYZTb+qIxHYYf2HlQ4fyxcV8B3
In8hSusO52CnHDuS+5w3YHMMDQDbj/aPztCz8hDf0NovyKz+g22bVW12xmMh
thydYT32JSKdKVNisRtC+pLtu2kSpgzEC7Ruxu/XTgfAgVsFCBeyKqqepbyI
2VIqtXCVDllFO24cd8Uxb549ACqAL1k6KKGEmlwV3K542aFkIWIuB8pKfE+P
BdWvokTmLP0C9pJVZdJ1YWbEMky+LoOwxS06bT2akYdBtijF83gWVwMEIYJo
hV3S4YHdqd0jv0BzwsUIoY9AdTC6v3vkCieYKO93VhzQ2fkdsduWh7vESEzs
VoIHL0Ser4baK1XOEfduW++WjHkcQpfYeRdR10FlagTF9M6m+/KdR5Koh8bv
fMDxBK5gV8k/ZkDH97nw+PTfYFhjw6u2BtpJMvYxfAj8BFUE0qGj16UDgSSk
vKo1GoWS2vxUVv2IkOZsiiYuCQsD6md0qtATtxovaobHNr2pnftS9Zt4Tzax
bk9bmfyMEbg02ddexLOJxk9BhsUc5zAATjQeXlA4giilj3j8mepK2GIWBr2x
x7sw8qXqNk/3h94etORxEMOc0Cj5hCNC8tCSi5aMQ9JPsHBsyzGkohwpj7/n
G7kWQpSHGvURxRLRTJSJZ0ub+aN8Yi41AMdxz1wcw/UX6YTKJcxpd3Z5SlI6
0p3zRyOjTqASsY7+8gjlvas4KkC6fuqrZKpn88zCC3b7oQ3s/7jMQx/m0MZa
FcUVYCRgAgiDipWRIFeDqjqeELfKzoy071HBbDbFsk2Ah62DMQIAww7bWKbf
9CGA7XNbxbtKnrxEoIlAOTAyLKJC7/MLiVro169qLaFJXqoJ9ssGXgpFS/df
ERuFcICiL/GFeXTvhHP7UDFK5dm4NmFeujcNXIUfLgOdso9cgBa4mxFfcAE4
d/MlJ+wEUS9WAQs4ZXSeL+sSXV050PwcnepM5aHBwJu4MiqELShiiPzKcKY4
w8JpVSISCVAQvnvLXRhFMrVsKJ026ETsO7yngHsodAL/1rfaD7YJb9Xj2L7A
4QknBLY3JP7EKbQHUrrYZXEZsZhrqXtkDOFOtL8faHpRwlF6Fcpbj/ai2bwK
Vsz6n5Hlv0Yovi/QI9rDHdBQ4EI4lPIOIKRx/NLFvAdx3U1W+rY7mpP+X0O0
OoS3RM7A4r1wYY6CRQvJwDV67hLnAAWCfMMq2cfLDzt77vPC3gM5o0bhmByU
/sWg+LpKE9GP6twL82J7EyY4iqH3Rq2GUvTcBzLBDF9H9iWTn46wuwbrLQXi
L54qs/U2/jaPt8rD7B2ilRFa5aRLv6JueyyVhTI2EG0eqMbepP6OZm1TDxCG
Zcj+rEyfwPXyxfeLIavDZ88eAL6ZQqbGb/GJfaQDEAElf6/vFzGO4ZSa/jc9
ziRlUZYlWjA6sNCCRle/ca2BIqGJh0w8dwsPWjOBgtdrl1IAY9BCymfjIfIS
Nzwu8AEVEKnU0lQ9+fiC4T7Njo8oLkShYK0+Z8p9PX94l4M4ldLmsjfIOsgv
y9db++Vk2WFeBDf/FTzOAjvcti0RjAYALufgVZTGsuF+61GD2OddSEl1mwT1
CBAwhr7eeDFURMaujZCZpYsOyQjDrCRbX70wQvIeOIBjtbksyvc4vbCnc59j
u2upgpCx8Ht/9OinO1Blebr37yiZwiNmaBprdwO0UzwRM26MovKy8DhjoDjr
NRH8hvSN5RB0ykWwOs6lfmLoADJE3PoKS5XqjwvpJYxijzyDYuN4fTGVeUin
RDY+85dozOcMAUzTnl9bG/TjBwpzyfIgR2hubCMI4TlLVgTStH6nS76TNKiR
xmi6pDbr7y6V9YfHkNqv++PnuFltfYuqoN35/nE5B+m9eNKshkBf+FoqWdve
+0S33IvUMrON7kxXIC8A4yGNSLtYcrRBcVwTt9ujNN/xuxkEO94HB8PepbOj
EhallxxwgbEZbXYnGSPfaoiOQuG4yIlnzUIJD/qYcEoyENHqq+RkkfJpF3cF
T586lsku1mYH22IhyMPvcxSUgY90KLKN8MwANJWDFZfWWAdIHOB35qQn4niF
itoARjMF5EGSvQIdwPAFMUeZtTyvPsVVLC4fWAnhWIPVn2L9XI3kxY+oOTri
8BPdXShAI9Yk/jRE2sTI+0T9b8YhlhVwkmtRXLXN6Vh03Q+HEObaXoMwSvhH
FDtqxn61zfNoxUY9UdQqYKiqaqMl5vOJlZnUSIoWKaFvVpnVRZhFXI51ouub
9FLkP/9oMf7B2gDr/BL3rvI3/lPGUSRDFK+7ApoHNMkYwqn4XJJkShqAsECv
2W7UEwdic3I4WC3zWPIqq7vkQ+AE5152gVCra9n2+chrOdYcwYbnykWPKo0Z
IbUFVnY4DPe+MCHK6YJpqoKdFFWgDkzeILYwGXjwwmdfL1x8YB6jYJRMHkpX
42yt/v6ZYmG9n6WZpW00pFZqy1K5uk3oMb7+xM4ZeDthFdDeLuw6Ql8QM3Dl
XDybvOij3GpGQEemLjVBr1vMfeNJJUlnIWp68nMEZbxtVtzY7FYRa9hdYw05
3q1MeLOWTNH6n4GpEdCRSXQEDDsqZLT4IG8AjO+Vdip3mdLojZCVeDkdLNIr
uxn764hxlPbWcXIAY0W8Iwbdb9Ri0eY7djBoJOfptCjKu8SggoUzXVrdqaUG
jVGZMAG0m+sruxYgwSKBgf0d2JlUKz8Mnf3FsCdTRFYHV5K/kMbkf9aqZA9m
LY48b9R/jFtXrR0xlW/9l7ycBunqmS5qxXNbxxMo/FZDrU8jOaxO157zolcv
7Eq+HA2r86QYjXAakKM8hX13sMM0fpzx8nxoCGRdrwiVAnoA7eSPjQrlz5Fz
VgoOKh2Sab++I0Nntl7LbYd+W65OStSjomd8+8ZmcyTgi/QthiJz4Tf7dEvW
tSdV/x8u9k9a80becr5Tv8CJocccmh+Nf+uD0pCfesaWkZMz6AkNV6BtmFFb
XmKcsTk28Pa5R7wRRHAKmZijRAS/+VOPTi2xnSeFXdEWfXutqPtGrTOBz7sg
E7q1J+L8w3pk9N3CxegGUzRgxj4IxTyF2+S/0kEdikLKOm1QmHlPbP3yP2no
KklanOkt3sCeLoFd+/ABt1sQFfgVDOS8/SzIrKiAUrQwh20adukGpdbXU8cB
KM3ryPT+2xDDJMiA0a77DGUMt4BI+LOzRf95aB7kZeIsxqJnS5cnsnBnCDzS
s/ohlVcj2DSYZ7jpgI9gV8ttpeB+aIUw4silun1ogXWdhY73RUt6x8b3JOfs
b8tcibFsJZy44u/Ntr3M+Ii7wu0xWEq59HzwOFA+UoJ12PpftBgvczArQq5m
WfFiYidYj008hczb2aBTpLEaGF5iszvUqymj7FvDJ6cLkrCk+gHc3PS/UX4W
HLwFNDmcjUb8wx2uVBnoWXbX8TzIFnHaqs4pg3ZveU1sVzLKsyiDyTvJbCHM
s8UjkHNST6rqxNFVxwSkHJDxSbCD9krKfHZS/t2pH/kFuNo4L3LjxaiLfkSL
rvbsCehf6tA+ObvhU7ObXrGNWY8lhJiaJEJvgpfqpmU9d+dX5+RBdmI+Stmr
mvytNRL1Ny4UUphkAWRZXQexsd/ZKnEkrzx8ws+xQ8U7R6R212tRTqJVRVG6
dgQTP1fiArMK0xbndbkOcz89LGcdPe1MymG0JsOyaA1j760YEeD+zaEUktI+
qHWIfIcdwKZh0MHbSPQ/UzdvcpqjMg/mQE/nWlYRIekVHh8vimnV+FyAFDux
Gd6l608lc7qs2g+pyROkZzZfy/I4LnqtawDWefU7CAMZTHpnj93TGbBWrkNV
OZzMPqmLXJM53QWNHJgWKapopMhbE/9WOPgUKx/HQVF8WDIle8xWXBsz9Rh8
LTmfdxn72b94PqntM3YPvxvT47HLRLQm6GCRgWBDGDZWHRDQ1hiik0C5yiuf
jKsQtmwHQL21iw5vjxHte7twSffrsbK9VTzBdqGgRxdbvVDvLxiK4u/dYwwu
BGHc3YGUlrTyGmFy55rmB8Mqcts1Pfv7j2OnKW7LSrjpIaW9Oj2B8DLsumgm
o745Nd0UAzo+zPmqKA1owVn0VgojTqxkJwGiR4MpiZMo/U01faC0gxsVfgJC
VznSeLkI7bjeZcHagNjXhNsT/aA9absjR98zU+J9k5wRzCKJ/MhZIkk+C3Ce
ZunQZKJqh77vWFwnL3L7SWtm6klmvkOTCjx0FDKHlnPZNvNw9+/1Iy7vM9nQ
Ps1kvdYhjest3IC4V6ZIV72pXYdvJnwXaL0TSGEX5NIQaqFC1BGI2A5KeZV5
7mY65iZjKPCS0xB4RZmHpxDR5cN28D4Bq5BnEj3Lr8Q2Ofqd3d4hNBWxT7hh
9KE5KgpdZlAFhk4K3ExBU1NeuW29v9q3U2+Ml2lyhDPwnNWI6djY4RkTsxNO
f7aZ2U96dZN94OKlEv0UuNE/AsS8CPAKOQ6sp5fzKp4dOgvRqtUtkh6fA1Fe
LEjKus4M9NYg36bAQQZjblC/al0BGrKFRlRf3wIpF1V7jDSZ24Et60ARNiPJ
4mtgQzLmo1V9CTSIa4xxIUBRQUjJ1sQw6bssojWP4gAqAZ4Ovqn691xWTc9t
Dd+tK9ww1e99lwir/7MkUpM2dR6JYyyRPLWu0W6ia/iPGznsqyKRyQebBNPh
MGjYjo15/MLgcc2wXd1A9B8msDiiYbZXVfJLZF8e7yw6vZC2iauKyAsznb9c
XkUln4fxS8/NhI5o4fnCmdlW8faR5sNgxHRdX002tmUUkuAPu3ucsNwt4qpn
+iurCnI2ADXWBgAAJwRhR479VnAUzqNEVOOMkaap/T0vLqFnke4NQxuigwKJ
ljhN3WIdq34rk0VM6e9nGFj+cTjHWQi9GKW7rqIfuKvSMIpo9RsfGbF7jyGf
xWMn2LcDz2VC3zsCS78SHB9cFNnk5wc4AKkckvEu0TYXWjAwfyv39kHlRb8s
xHkVg0sjWieQOYff7AkMAwq0QqHmO2F0r/E+vGbzZkrvYZBXjLhNICF5zeRL
GjRfo4+PRLAZNENK2P3rIw/z10VBY09PpnTftfpy04Muf59UHFlRZzcSa8Mp
BD+CAjguO28kFtJowCPsyjb9IjAtmvigT7BceZwiQgXqZMTm2tVbhrkKpkdw
QGbKhUJvlpenejlAMc6BYETQc9BIlVgJYA83aKwdAYnoa21CTKagTrmYms5S
IEfp5bsADNNEIyHYpbcXKZivhKCrX3K/Qlx+AN6gDHhac6IhL0sY7R8vTjkK
eA+mhYZJqIaYvY9ZG0FSkCJf7Ib4o4qBhOJq8WQ3WL9bg86eUbG8kYWnLjE/
Ul1K6jg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe76PxC8qxyheZ1lwMfdUwSB7bsYZt16f0THHoKZq2AwxQkDdhDzG4hPIkahiOMFgv69TmWdKMATMtc9eNHzAYxwp28dgkSzHQlzxufI99CsatB5/IcJekwRRYokLCL3qmjxEc7vPUeeVRrwJQwlySvSXNqL5ytpM6uOE1UIbyGoo0KqC3wuyoIsQTMlerIdcvKa2b1DM1m3R/jrLC7ObscCXFnxuRD1blnBKj9QxUuCzPfshCVf2aoKgSFZ3i51Q0OZVZfdihipNYEDIMd8z9d3ZAINI8OV1rdZQ/QXtJ8zNTciXUgIMculfCLQJk7GCl8Ey8dR+7RBgllb4SnCf/OGoKGnU5amnPMPOw5tYBRXR7I0S3GWkF90I2fzBFLe0davR/bIZ7fORA8RUNzq8F9gQ5dZpwy5+PN3BQch6pw5RP2JBUEbfC7ULCTRstiV21fwUkfjAjop6NqsgnrRCTprKZJ2q8e4oCzb6BiP4O/BfYXgdnoIRruCXHsXEun0sWz9TKHfv6l9N981A+sCmOBtKySgKdsJHdTC96jtdCr5pSnr/35CQ/LK91vdVoYy0ATM8J5wK10arUr8QFcwuoyCe6TG3BnmXnseKyTb0a8SflfVK5on0EYMUQsMLbPnuC4M3FMq7yX3S/iaQf7YV0I1o+BvAE5BpXUI6LBRRKm83XmRmXk490evlDsXbBdyU+Na/XjBdIeF2+9Lq5t5Y444MDs2ZgoruatPRHKHNL5gRAAcW8Urs36vEQ9/RrkuBYB8y7LcvmvVvlkVo8H9Huoe9"
`endif
//########################################################################
//# Copyright (C) 2025 Altera Corporation.
//# SPDX-License-Identifier: MIT
//#########################################################################

// `define SVT_AXI_MAX_NUM_MASTERS_1
// `define SVT_AXI_MAX_NUM_SLAVES_1
// 
// `define SVT_AXI_MAX_ADDR_WIDTH 64
// 
// `define SVT_AXI_MAX_DATA_WIDTH 256

`define SVT_AXI_WSTRB_WIDTH 16

`define SVT_AXI_MAX_BURST_LENGTH_WIDTH 10

`ifndef SM_ETH_AXI_SYS_SEQUENCER
  `define SM_ETH_AXI_SYS_SEQUENCER env.axi_system_env.sequencer
`endif

`ifndef SM_ETH_AXI_MST_SEQUENCER
  `define SM_ETH_AXI_MST_SEQUENCER axi_system_env.master[0].sequencer
`endif

`ifndef SM_ETH_AXI_SLV_SEQUENCER
  `define SM_ETH_AXI_SLV_SEQUENCER axi_system_env.slave[0].sequencer
`endif

`ifndef SM_ETH_QSYS_TOP
  `define SM_ETH_QSYS_TOP tb_top.dut.soc_inst
`endif

`ifndef SM_ETH_QSYS_TOP_MM_INT_SS_F2H_AXI4
  `define SM_ETH_QSYS_TOP_MM_INT_SS_F2H_AXI4(sig) `SM_ETH_QSYS_TOP.mm_interconnect_2_subsys_hps_f2sdram_adapter_axi4_sub_``sig``
`endif

`ifndef SM_ETH_DUT_IOPLL
  `define SM_ETH_DUT_IOPLL `SM_ETH_QSYS_TOP.iopll_0
`endif

`ifndef SM_ETH_SSGDMA_PATH
  `define SM_ETH_SSGDMA_PATH `SM_ETH_QSYS_TOP.subsys_ssgdma.ssgdma
`endif

`ifndef SM_ETH_HSSI_SS0_PATH
  `define SM_ETH_HSSI_SS0_PATH tb_top.dut.gen_mulit_inst[0].hssi_ss_top
`endif

`ifndef SM_ETH_MOD_DEVKIT
`ifndef SM_ETH_HSSI_SS1_PATH
  `define SM_ETH_HSSI_SS1_PATH tb_top.dut.gen_mulit_inst[1].hssi_ss_top
`endif
`endif

`ifndef SM_ETH_EHIP_PORT0
  `define SM_ETH_EHIP_PORT0 `SM_ETH_HSSI_SS0_PATH.u0
`endif

`ifndef SM_ETH_EHIP_PORT1
  `define SM_ETH_EHIP_PORT1 `SM_ETH_HSSI_SS1_PATH.u0
`endif

`ifndef SM_ETH_F2H_CLK
  `define SM_ETH_F2H_CLK dut.clk_bdg_100_clk
`endif

`ifndef SM_ETH_H2F_CLK
  `define SM_ETH_H2F_CLK dut.clk_bdg_125_clk
`endif

`ifndef NUM_D2H_ST_PORTS
  `define NUM_D2H_ST_PORTS 1
`endif

`ifndef NUM_H2D_ST_PORTS
  `define NUM_H2D_ST_PORTS 1
`endif

`ifndef SM_ETH_SFP_DUT_PATH
  `define SM_ETH_SFP_DUT_PATH tb_top.dut.sfp_top_inst
`endif

// ------------------------------- CSR ---------------------------------------
`ifndef SM_ETH_SSGDMA_CSR_ADDR
  `define SM_ETH_SSGDMA_CSR_ADDR 'h4500_0000
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_ADDR
  `define SM_ETH_SSGDMA_CSR_D2H0_ADDR 'h4520_0000
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_ADDR
  `define SM_ETH_SSGDMA_CSR_D2H1_ADDR 'h4520_0800
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_ADDR
  `define SM_ETH_SSGDMA_CSR_H2D0_ADDR 'h4524_0000
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_ADDR
  `define SM_ETH_SSGDMA_CSR_H2D1_ADDR 'h4524_0800
`endif

// Device port CSR offsets
// addr [10:0]  register offset for ports
// addr [14:11] port number
// addr [17:15] reserved
// addr [19:18] 0 - d2h st, 1 h2d st

// ------------------------- D2H0 --------------------------------------------
`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_START_ADDR_L
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_START_ADDR_L (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h8)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_START_ADDR_H
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_START_ADDR_H (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'hC)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_SIZE
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_SIZE (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h10)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_INSERT_POINTER
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_INSERT_POINTER (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h18)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_RESP_SIZE
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_RESP_SIZE (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h3C)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_RESPONDER_ADDR_L
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_RESPONDER_ADDR_L (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h400)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_RESPONDER_ADDR_H
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_RESPONDER_ADDR_H (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h404)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_CTRL
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_CTRL (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h0)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H0_Q_STATUS
  `define SM_ETH_SSGDMA_CSR_D2H0_Q_STATUS (`SM_ETH_SSGDMA_CSR_D2H0_ADDR + 'h4)
`endif

// ------------------------- H2D0 --------------------------------------------
`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_START_ADDR_L
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_START_ADDR_L (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h8)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_START_ADDR_H
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_START_ADDR_H (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'hC)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_SIZE
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_SIZE (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h10)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_INSERT_POINTER
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_INSERT_POINTER (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h18)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_RESP_SIZE
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_RESP_SIZE (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h3C)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_RESPONDER_ADDR_L
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_RESPONDER_ADDR_L (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h400)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_RESPONDER_ADDR_H
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_RESPONDER_ADDR_H (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h404)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_CTRL
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_CTRL (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h0)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D0_Q_STATUS
  `define SM_ETH_SSGDMA_CSR_H2D0_Q_STATUS (`SM_ETH_SSGDMA_CSR_H2D0_ADDR + 'h4)
`endif

// ------------------------- D2H1 --------------------------------------------
`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_START_ADDR_L
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_START_ADDR_L (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h8)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_START_ADDR_H
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_START_ADDR_H (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'hC)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_SIZE
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_SIZE (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h10)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_INSERT_POINTER
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_INSERT_POINTER (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h18)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_RESP_SIZE
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_RESP_SIZE (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h3C)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_RESPONDER_ADDR_L
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_RESPONDER_ADDR_L (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h400)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_RESPONDER_ADDR_H
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_RESPONDER_ADDR_H (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h404)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_CTRL
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_CTRL (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h0)
`endif

`ifndef SM_ETH_SSGDMA_CSR_D2H1_Q_STATUS
  `define SM_ETH_SSGDMA_CSR_D2H1_Q_STATUS (`SM_ETH_SSGDMA_CSR_D2H1_ADDR + 'h4)
`endif

// ------------------------- H2D1 --------------------------------------------
`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_START_ADDR_L
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_START_ADDR_L (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h8)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_START_ADDR_H
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_START_ADDR_H (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'hC)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_SIZE
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_SIZE (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h10)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_INSERT_POINTER
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_INSERT_POINTER (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h18)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_RESP_SIZE
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_RESP_SIZE (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h3C)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_RESPONDER_ADDR_L
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_RESPONDER_ADDR_L (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h400)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_RESPONDER_ADDR_H
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_RESPONDER_ADDR_H (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h404)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_CTRL
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_CTRL (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h0)
`endif

`ifndef SM_ETH_SSGDMA_CSR_H2D1_Q_STATUS
  `define SM_ETH_SSGDMA_CSR_H2D1_Q_STATUS (`SM_ETH_SSGDMA_CSR_H2D1_ADDR + 'h4)
`endif

// ---------------------------------------------------------------------------
`ifndef SM_ETH_SSGDMA_CSR_CTRL
  `define SM_ETH_SSGDMA_CSR_CTRL (`SM_ETH_SSGDMA_CSR_ADDR + 'h100)
`endif

`ifndef SM_ETH_SSGDMA_CSR_IP_PARAM
  `define SM_ETH_SSGDMA_CSR_IP_PARAM (`SM_ETH_SSGDMA_CSR_ADDR + 'h11C)
`endif

`ifndef SM_ETH_DMA_H2D0_DA
  `define SM_ETH_DMA_H2D0_DA 'h0011_2233
`endif

`ifndef SM_ETH_DMA_H2D0_SA
  `define SM_ETH_DMA_H2D0_SA 'h0022_3344
`endif

`ifndef SM_ETH_DMA_H2D1_DA
  `define SM_ETH_DMA_H2D1_DA 'h1111_2233
`endif

`ifndef SM_ETH_DMA_H2D1_SA
  `define SM_ETH_DMA_H2D1_SA 'h1122_3344
`endif

`ifndef SM_ETH_DMA_D2H0_DA
  `define SM_ETH_DMA_D2H0_DA 'h1122_2233
`endif

`ifndef SM_ETH_DMA_D2H0_SA
  `define SM_ETH_DMA_D2H0_SA 'h1133_3344
`endif

`ifndef SM_ETH_DMA_D2H1_DA
  `define SM_ETH_DMA_D2H1_DA 'h2211_2233
`endif

`ifndef SM_ETH_DMA_D2H1_SA
  `define SM_ETH_DMA_D2H1_SA 'h2222_3344
`endif

`ifndef SM_ETH_TYPE
  `define SM_ETH_TYPE 'h800
`endif

// ---------------------------------------------------------------------------
`define MULTI_EOP_SOP

// --------HSSI---------------------------------------------------------------
`ifndef SM_ETH_HSSI_CSR_PORT0_SOFT_IP_BASE
  `define SM_ETH_HSSI_CSR_PORT0_SOFT_IP_BASE 'h4030_0100
`endif

`ifndef SM_ETH_HSSI_CSR_PORT0_HARD_IP
  `define SM_ETH_HSSI_CSR_PORT0_HARD_IP 'h4032_0000
`endif

`ifndef SM_ETH_HSSI_CSR_PORT0_HARD_IP_EMAC
  `define SM_ETH_HSSI_CSR_PORT0_HARD_IP_EMAC 'h4035_0000
`endif

`ifndef SM_ETH_HSSI_CSR_PORT1_SOFT_IP_BASE
  `define SM_ETH_HSSI_CSR_PORT1_SOFT_IP_BASE 'h4050_0100
`endif

`ifndef SM_ETH_HSSI_CSR_PORT1_HARD_IP
  `define SM_ETH_HSSI_CSR_PORT1_HARD_IP 'h4052_0000
`endif

`ifndef SM_ETH_HSSI_CSR_PORT1_HARD_IP_EMAC
  `define SM_ETH_HSSI_CSR_PORT1_HARD_IP_EMAC 'h4055_0000
`endif

// --------ETH BRIDGE / PKT CLIENT--------------------------------------------
`ifndef SM_ETH_BRIDGE_CSR_BASE
  `define SM_ETH_BRIDGE_CSR_BASE 'h5001_0000
`endif

`ifndef SM_ETH_BRIDGE_TCAM0_CSR_BASE
  `define SM_ETH_BRIDGE_TCAM0_CSR_BASE (`SM_ETH_BRIDGE_CSR_BASE + 'h100)
`endif

`ifndef SM_ETH_BRIDGE_TCAM0_CSR_LAST_ADDR
  `define SM_ETH_BRIDGE_TCAM0_CSR_LAST_ADDR (`SM_ETH_BRIDGE_CSR_BASE + 'h40FC)
`endif

`ifndef SM_ETH_BRIDGE_TCAM0_KEY_CSR_ADDR
 `define SM_ETH_BRIDGE_TCAM0_KEY_CSR_ADDR (`SM_ETH_BRIDGE_TCAM0_CSR_BASE+'h1000)
`endif

`ifndef SM_ETH_BRIDGE_TCAM0_RESULT_CSR_ADDR
 `define SM_ETH_BRIDGE_TCAM0_RESULT_CSR_ADDR (`SM_ETH_BRIDGE_TCAM0_CSR_BASE+'h2000)
`endif

`ifndef SM_ETH_BRIDGE_TCAM0_MASK_CSR_ADDR
 `define SM_ETH_BRIDGE_TCAM0_MASK_CSR_ADDR (`SM_ETH_BRIDGE_TCAM0_CSR_BASE+'h3000)
`endif

`ifndef SM_ETH_BRIDGE_TCAM1_CSR_BASE
  `define SM_ETH_BRIDGE_TCAM1_CSR_BASE (`SM_ETH_BRIDGE_CSR_BASE + 'h4200)
`endif

`ifndef SM_ETH_BRIDGE_TCAM1_CSR_LAST_ADDR
  `define SM_ETH_BRIDGE_TCAM1_CSR_LAST_ADDR (`SM_ETH_BRIDGE_CSR_BASE + 'h81FC)
`endif

`ifndef SM_ETH_BRIDGE_TCAM1_KEY_CSR_ADDR
 `define SM_ETH_BRIDGE_TCAM1_KEY_CSR_ADDR (`SM_ETH_BRIDGE_TCAM1_CSR_BASE+'h1000)
`endif

`ifndef SM_ETH_BRIDGE_TCAM1_RESULT_CSR_ADDR
 `define SM_ETH_BRIDGE_TCAM1_RESULT_CSR_ADDR (`SM_ETH_BRIDGE_TCAM1_CSR_BASE+'h2000)
`endif

`ifndef SM_ETH_BRIDGE_TCAM1_MASK_CSR_ADDR
 `define SM_ETH_BRIDGE_TCAM1_MASK_CSR_ADDR (`SM_ETH_BRIDGE_TCAM1_CSR_BASE+'h3000)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_CSR_BASE
  `define SM_ETH_PKT_CLIENT_0_CSR_BASE 'h5000_0000
`endif

`ifndef SM_ETH_PKTCLI0_CFG_PKT_CL_CTRL
  `define SM_ETH_PKTCLI0_CFG_PKT_CL_CTRL (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h00)
`endif

`ifndef SM_ETH_PKTCLI0_DYN_DMAC_ADDR_U
 `define SM_ETH_PKTCLI0_DYN_DMAC_ADDR_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h0C)
`endif

`ifndef SM_ETH_PKTCLI0_DYN_DMAC_ADDR_L
 `define SM_ETH_PKTCLI0_DYN_DMAC_ADDR_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h10)
`endif

`ifndef SM_ETH_PKTCLI0_DYN_SMAC_ADDR_U
 `define SM_ETH_PKTCLI0_DYN_SMAC_ADDR_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h14)
`endif

`ifndef SM_ETH_PKTCLI0_DYN_SMAC_ADDR_L
 `define SM_ETH_PKTCLI0_DYN_SMAC_ADDR_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h18)
`endif

`ifndef SM_ETH_PKTCLI0_DYN_PKT_NUM
 `define SM_ETH_PKTCLI0_DYN_PKT_NUM (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h1C)
`endif

`ifndef SM_ETH_PKTCLI0_DYN_PKT_SIZE_CFG
 `define SM_ETH_PKTCLI0_DYN_PKT_SIZE_CFG (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h20)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_TX_SOP_CNT_L
  `define SM_ETH_PKTCLI0_STAT_TX_SOP_CNT_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h24)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_TX_SOP_CNT_U
  `define SM_ETH_PKTCLI0_STAT_TX_SOP_CNT_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h28)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_TX_EOP_CNT_L
  `define SM_ETH_PKTCLI0_STAT_TX_EOP_CNT_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h2C)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_TX_EOP_CNT_U
  `define SM_ETH_PKTCLI0_STAT_TX_EOP_CNT_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h30)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_RX_SOP_CNT_L
  `define SM_ETH_PKTCLI0_STAT_RX_SOP_CNT_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h3C)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_RX_SOP_CNT_U
  `define SM_ETH_PKTCLI0_STAT_RX_SOP_CNT_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h40)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_RX_EOP_CNT_L
  `define SM_ETH_PKTCLI0_STAT_RX_EOP_CNT_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h44)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_RX_EOP_CNT_U
  `define SM_ETH_PKTCLI0_STAT_RX_EOP_CNT_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h48)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_CHK_MISC
  `define SM_ETH_PKTCLI0_STAT_CHK_MISC (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h58)
`endif

`ifndef SM_ETH_PKTCLI0_STAT_CHK_CNT
  `define SM_ETH_PKTCLI0_STAT_CHK_CNT (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h5c)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_RX_BYTE_CNT_L
  `define SM_ETH_PKT_CLIENT_0_RX_BYTE_CNT_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h60)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_RX_BYTE_CNT_U
  `define SM_ETH_PKT_CLIENT_0_RX_BYTE_CNT_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h64)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_TX_BYTE_CNT_L
  `define SM_ETH_PKT_CLIENT_0_TX_BYTE_CNT_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h68)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_TX_BYTE_CNT_U
  `define SM_ETH_PKT_CLIENT_0_TX_BYTE_CNT_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h6C)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_TX_NUM_TICKS_L
  `define SM_ETH_PKT_CLIENT_0_TX_NUM_TICKS_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h70)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_TX_NUM_TICKS_U
  `define SM_ETH_PKT_CLIENT_0_TX_NUM_TICKS_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h74)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_RX_NUM_TICKS_L
  `define SM_ETH_PKT_CLIENT_0_RX_NUM_TICKS_L (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h78)
`endif

`ifndef SM_ETH_PKT_CLIENT_0_RX_NUM_TICKS_U
  `define SM_ETH_PKT_CLIENT_0_RX_NUM_TICKS_U (`SM_ETH_PKT_CLIENT_0_CSR_BASE+'h7C)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_CSR_BASE
  `define SM_ETH_PKT_CLIENT_1_CSR_BASE 'h5000_1000
`endif

`ifndef SM_ETH_PKTCLI1_CFG_PKT_CL_CTRL
 `define SM_ETH_PKTCLI1_CFG_PKT_CL_CTRL (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h00)
`endif

`ifndef SM_ETH_PKTCLI1_DYN_DMAC_ADDR_U
 `define SM_ETH_PKTCLI1_DYN_DMAC_ADDR_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h0C)
`endif

`ifndef SM_ETH_PKTCLI1_DYN_DMAC_ADDR_L
 `define SM_ETH_PKTCLI1_DYN_DMAC_ADDR_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h10)
`endif

`ifndef SM_ETH_PKTCLI1_DYN_SMAC_ADDR_U
 `define SM_ETH_PKTCLI1_DYN_SMAC_ADDR_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h14)
`endif

`ifndef SM_ETH_PKTCLI1_DYN_SMAC_ADDR_L
 `define SM_ETH_PKTCLI1_DYN_SMAC_ADDR_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h18)
`endif

`ifndef SM_ETH_PKTCLI1_DYN_PKT_NUM
 `define SM_ETH_PKTCLI1_DYN_PKT_NUM (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h1C)
`endif

`ifndef SM_ETH_PKTCLI1_DYN_PKT_SIZE_CFG
 `define SM_ETH_PKTCLI1_DYN_PKT_SIZE_CFG (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h20)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_TX_SOP_CNT_L
  `define SM_ETH_PKTCLI1_STAT_TX_SOP_CNT_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h24)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_TX_SOP_CNT_U
  `define SM_ETH_PKTCLI1_STAT_TX_SOP_CNT_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h28)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_TX_EOP_CNT_L
  `define SM_ETH_PKTCLI1_STAT_TX_EOP_CNT_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h2C)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_TX_EOP_CNT_U
  `define SM_ETH_PKTCLI1_STAT_TX_EOP_CNT_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h30)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_RX_SOP_CNT_L
  `define SM_ETH_PKTCLI1_STAT_RX_SOP_CNT_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h3C)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_RX_SOP_CNT_U
  `define SM_ETH_PKTCLI1_STAT_RX_SOP_CNT_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h40)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_RX_EOP_CNT_L
  `define SM_ETH_PKTCLI1_STAT_RX_EOP_CNT_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h44)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_RX_EOP_CNT_U
  `define SM_ETH_PKTCLI1_STAT_RX_EOP_CNT_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h48)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_CHK_MISC
  `define SM_ETH_PKTCLI1_STAT_CHK_MISC (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h58)
`endif

`ifndef SM_ETH_PKTCLI1_STAT_CHK_CNT
  `define SM_ETH_PKTCLI1_STAT_CHK_CNT (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h5c)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_RX_BYTE_CNT_L
  `define SM_ETH_PKT_CLIENT_1_RX_BYTE_CNT_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h60)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_RX_BYTE_CNT_U
  `define SM_ETH_PKT_CLIENT_1_RX_BYTE_CNT_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h64)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_TX_BYTE_CNT_L
  `define SM_ETH_PKT_CLIENT_1_TX_BYTE_CNT_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h68)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_TX_BYTE_CNT_U
  `define SM_ETH_PKT_CLIENT_1_TX_BYTE_CNT_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h6C)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_TX_NUM_TICKS_L
  `define SM_ETH_PKT_CLIENT_1_TX_NUM_TICKS_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h70)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_TX_NUM_TICKS_U
  `define SM_ETH_PKT_CLIENT_1_TX_NUM_TICKS_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h74)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_RX_NUM_TICKS_L
  `define SM_ETH_PKT_CLIENT_1_RX_NUM_TICKS_L (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h78)
`endif

`ifndef SM_ETH_PKT_CLIENT_1_RX_NUM_TICKS_U
  `define SM_ETH_PKT_CLIENT_1_RX_NUM_TICKS_U (`SM_ETH_PKT_CLIENT_1_CSR_BASE+'h7C)
`endif
// --------PTP BRIDGE / PKT CLIENT--------------------------------------------

// --------USER SPACE CSR--------------------------------------------
`ifndef SM_ETH_USER_CSR
  `define SM_ETH_USER_CSR  'h4020_0000
`endif

`ifndef SM_ETH_USER_CSR_CTRL_REG
  `define SM_ETH_USER_CSR_CTRL_REG `SM_ETH_USER_CSR
`endif

`ifndef SM_ETH_USER_CSR_ERROR_REG
  `define SM_ETH_USER_CSR_ERROR_REG (`SM_ETH_USER_CSR+'h4)
`endif

`ifndef SM_ETH_USER_CSR_STATUS_REG
  `define SM_ETH_USER_CSR_STATUS_REG (`SM_ETH_USER_CSR+'h8)
`endif
// --------USER SPACE CSR--------------------------------------------

//------------------------SFP/SFP-----------------------------//
`ifndef SM_ETH_SFP_SYSTEM_OFFSET
  `define SM_ETH_SFP_SYSTEM_OFFSET 'h4404_0000
`endif

`ifndef SM_ETH_SFP_CFG_REG
  `define SM_ETH_SFP_CFG_REG (`SM_ETH_SFP_SYSTEM_OFFSET + 'h20)
`endif

`ifndef SM_ETH_SFP_TFR_CMD
  `define SM_ETH_SFP_TFR_CMD (`SM_ETH_SFP_SYSTEM_OFFSET + 'h40)
`endif

`ifndef SM_MSGDMA_DESCR_LENGTH
  `define SM_MSGDMA_DESCR_LENGTH 512
`endif

`ifndef SM_MSGDMA_NUM_OF_PORTS
  `define SM_MSGDMA_NUM_OF_PORTS 1
`endif

//------------------------SFP/SFP-----------------------------//

// dma addressing: 31: 0; [30:28]: DESCR/DMA_DATA; [27:26]: H2D/D2H
//                 [25:22]: PORT#; [21:0]: $
`define D2H_ST_AGENT 2'd0
`define H2D_ST_AGENT 2'd1

`define DESCR	   3'd1
`define DMA_DATA 3'd2
`define RESP     3'd3

parameter PORT0_TXDMA_ADDR 			= 32'h2400_0000;
parameter PORT0_RXDMA_ADDR 			= 32'h2000_0000;
parameter PORT0_SA				= 48'hAAAA_AAAA_AAAA;
parameter PORT0_DA				= 48'hDDDD_DDDD_DDDD;
parameter PORT0_START_DESC_CTRL		= 32'hC000_1300;
parameter PORT0_END_DESC_CTRL			= 32'h8000_1300;
parameter DMA_PORT0_BASE_TXDMA_PREF_ADDR       = 64'h448_0000;
parameter DMA_PORT0_BASE_TXDMA_CSR_ADDR        = 64'h448_0020;
parameter DMA_PORT0_BASE_RXDMA_PREF_ADDR       = 64'h448_0080;
parameter DMA_PORT0_BASE_RXDMA_CSR_ADDR        = 64'h448_00A0;
parameter DMA_PORT0_BASE_ADDR       = 64'h448_0000;
parameter PORT0_TXDESC_BASE_ADDR      = 64'h1400_0000;
parameter PORT0_RXDESC_BASE_ADDR      = 64'h1000_0000;

//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OPyG3vzrwPsOWGItA0ia8DOJfkWt7W3yj1Qkhkz+ykPTphYM8ypPS5MPFrxT
Jb76LU1O/H+ABhxyeUGd5QUhdQsCG8dzVRQkhOIJDhCfWWW1IOm/BVqaSzV+
+YAkQSzT8UaE12+WYhvBEOdpfcZ7Q11t1URr6xec/gmt5L2vDDjtmv7kEeRw
LAaH96MD44ygAAmE46lqQDzxVOM/vbU7s0VWo8OR3aZSfp80dv9cw9PKiFaR
uT4taP/sTj+PI3rJo44gKH+cAlOqnIdPusH6C3E/G1wjEn0pqgFXUWSPtPlT
wl1qKeiD1fgrD/5umhltSMPMuU9JQk735GgWsyamwg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FWtBHqCAjXm+QUxHBHJc1qQePPGoE8NQmryoTyek4/d58mDQ5cxjiOd2p/HH
lEKOUYLkE342VIFW6q9wuHITBRGLcHEMOrpl/e82LDJLQsAY1FwtiBamQiCB
vxu2JwnaFQXH6NoNV1msDrnYpJTuYPveD3TGsOokYpmSYsGdpI48XrewM/1l
24GEp5cN9uP1GG0unxO78OCzWif18wLeKEjM/Fe1xurKPPmfcBFTYEEIg+R1
JcmQwnDBmRQmLK4yg6ScAN8pgNwZbJEUfH8WtW65tAGqAkLsihqHzfR53WSZ
M5iV7Tn5cgjXVHbFkoTUC2hqDFKvQMqMqJSFNTZpgA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I2hkDfYQqrTrEg6GA/vzRFfY+Tg4ZmvmFlNNygBDui6SyhwVgoEOJl15l/7b
zjBSfYUfoFGILtulMWcdJcfbE4MKRhy4Ho5iPEVqkTvx+VZrLlvNWC3XmXZM
2pXkb+cyJHxWCeIvzZ3pxBbSz56p/zM1WihYbKTEPI++JVLH3o26GdXmO0/b
zV1yRawUvRuHRitO5440pr4CCjCnzUCMrj+BmI+XVwapq8uEhG7GwSZazZ6X
WlPetXds8ClqbJh4PBLGg7IH9skkajQGp71hOwDo2hUD1CrjYtUiO5hKVT8v
ifEqk5DdeuZYGxFiWpFrf2dEIZa123WYkTZ93Qbd1A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mXecucQjarMhBnLDJudlCjW/vuMeLGiuPUdPhh1MKFoKilIV/h/tdpLZP0nV
rJkm0RZMBDt+hOqipHDAF14dwOg6ksXua1cCef84NhxQHafy3PQpx/tGQQlb
6XYkbwCpUlbhcq07eckfNHHFDJmARLt8QRmEzdnoFsMiLfLnz1xzbyY/ydf1
9oyFsTu7HwBxux1TYbJfx6wef/6IgEOBE/xYwUfzFlyBAJr4xPWL55ZVKrbX
hGjNO7DI+t3uNqxXrRvdaCFznaQ0CTeDR45x0SC3rehZaSq4SgZIr3ohbZJ1
2qy3NRp4w1VvO2wCawsP4vaOytPvAJvxqG51MBi9Ng==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZqvM1Hm73cODASMa1zQWby6UYw+J68tm5htUpMBr9G7wQLD5nNWyYYgdgkTL
FM6d/LWeB0FDQlY6ZPE2xP7wYwnDhTBr5Be6CaFJV6fIlriLzryhnvMY3O/U
ksuMgHswYuT+dSjsZgOqvM1K+Jay3Nm6+P5tR4+bYd2cJ+Jn6ck=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
fOr7ReNKclhM8qumBzeAoLz6hhg2KV3i/9qOgxyIAETPIPa2y7qUGGebEYcx
Q6FrrD0FqEHItlwaEc2y0m+EJ4aaLy4OFuqgKmwCH/YcWjdsbb8it6ja2Tby
cQnrJkr1JSg/APqnHCXDywERrTGwGxzkkfyQxWMUtbloLvYgiysOTCzSdXgp
ojMXUEo+Di4wfUpO9aBlaD9dhLunotnuFtjRNiO5fhVe+Q6KnDodMOWuY/UF
lfOzGUoClQRSuaQMPLvwF/1WGEdlyVtE8X1yzLtb956rdTJRcMs1XXUdn8FL
0paRk3zzeTtXGPGmxrDI885iE9rr0KHtTaA/NyS8LGrtApgX138ReLCRHz9C
uNsqGa6zK0yxOJE7/TosZlUhtiu0sZ6X3u2nKxQLeCFK29nskGaf0RMoblos
8wmnazi7XHr5D+xnTxQAhSh4jXyjNEFxeAZILiIfAj0qDeKJ9gSS/Sg7Ky8T
xQ3juA+bX3mdMbIMOcbXZ7ss+A06HJXU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BlnYi3wagmCOudx6Lw+3Y1HVnU1pUBYE/Q2KplxXYLDyp3KLRXTyRv7pa3LI
etNTSm3nakqIhG4jj4iIMLfIAvdq54EvtyOm6m1+ZFuigZ9lJ7+j21xfHBQY
q26Jvaq+tIgWlNdhe/PWxKUeMjoWEj7Y4vT4m1cT2A6ay1Uz57Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FDWfG+jmF/MatBudEJeGejCmXuh9B2P34aVWgqSlGOUjo2bz+M9BRslpR+B/
tq0LwjbIQDO2KNPzy4kaZDVAfvYChupfy4picUsgCjEV049Yuq761XhNVq0L
0qNAftcrKHQOlzYy4xnrML1OswmOLqU2H1rLJLb0FfBefUG/LPc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
lPmsCzsAo5uGbdJGitv0j5ayJny7t5xcVryBpuorEU4kLIvpCS07GLKIIhz+
TRiPzfXpCdJ3trRKPKmhFL9wAr8gtC0uO0G5stp62AN5iDZb7V+d53bUTW5W
6oVYdhWKosgA28IEJAxCIGAQYHwnqP/YHm5Nl37FImxBBVRGPBiONWa1WMMd
wewcLfhQdiIGH5QeEMciII7MCQFcCE4kuj3nIA5Y9uADwYijwfRoUcFWQWtq
oDDjLmaDpI3gH6mhEVK5lSViNI2np0a+APQt/IFXpe/bd/+fzRE47WkZUmWa
dLiasYTKg1+j8WOSmOXfWNNV0pPeetiGczDfQ6k1fl52hi1NH2Hsgym3ZMPf
tkyOwYkdCj9O1rpZlEgHl4W3QZrFqzOIw5eY2DBzcqZWIBOO7wEaRYbobunC
TMdsLTERRGUziVqHXJ52davdQTF0DHgVvIeoSk7DqD6aGUs1W8fWucPwinXP
l7mOLLYha6LTVvX5EMIbNRn2yxmq9KeACSNj+OzaU3Mfr8G1cPtxGiUBtm9Y
w7EInFVd1prtFPDpfc4leNiif4ZCv75FGiEpTScB2UchCfwkLA9pLJ0wfUyO
Gqojv9IrKiY25/Zp0pxm25lOBaWopaKfrWQ4QSj+vqDkegYeOWGb5USIbs28
eCCOxxcBCM1UkMidC75RbbJKRMayp3xc9rRtzRvnBq87LqyznZNHVHDWVKQJ
WA7TV+zXsZHDH+BVJd9Vo+BJg6d8MPfdgMRMWQ7BGkpYG1AJaOBUgNpuy2ea
fdr2MvSNPZhgr0a9J3y+kQcFEOuU365ECmv/XG6PfDdpFAA4BITuJ8stl3y4
7swc48APx7yWzzdj4Ss5G+JgCU/6/Be4K1deyu6nimta2ogoIzDwM92Tn/XM
fUgKGrjClwbfUTabN2/6paCxo3xKbu7/lzYyuRzqKFpi/UduOlxHdsy8yCZz
tYm1rCvwdVqkijuqKulzbcjXICqvueIIOAjCrD3iCQlXLDi8bvDHHxFI829I
sjSRqHAnz9jzy4/YsRDIPqikMq38wPoRMC6xhvRPn7ihIA4fZZifPAsyCOZ9
WRr7yZFWutJt9Ro1CpaVxAVbYhh8cHjFrn+j7QIRQzkJUgBZ/wnIC3c18qif
n9n3g7CcCZ9vgGj0NkGrhrX4a5/dDQ74FMObuK1x1f3SJNzcKe+UFr5rBtAy
31JmIcMU1udNa7ucfk3MVwlaMu8GHabwoucSER2/K4XEOGLclk4hSRL6MUep
mgVrReZU7XBtJuAAFkAtyy+wbxJVKriF5TeF0IaK3Yu0Edqduu+w/T8h750R
UK+QyzEB/xNCyX4cU0C8iW5K9eI892+ykzsDiDAQoLL94/8bHuI98D98sDZq
YavYJiiJvdgWOsyBBiVAPZ/3pliONjyhnlc1qVyE5g/VsR38ha8NVtpPIkjk
IDBYtmtBcFb8C1EMf3yeYHFN7FgLod17OyLxx9mVvq0FLBP/so4ZV1bSRncO
QOo0g0Mk12swy0H/Sc8AHULbPLgPRpaBn+oxAmUR9XbbQsRGjaCR3mKJ7eDK
hp8egtV6MZQxmoS9Xwd4xop5u+PaM221C7r1qjW0pd28NM2139aX4F58bzgb
auAbj4rIzPQeEUsNj+vyQIgnGOiQgrWqlgLi93UDljj1/+7uDDJ0fqd9eiwx
venAzGRZN073wKSBAblB1nzMMo4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe75bgRW2M6DGSLf3/XovlHu8yjibi20I2Vkq938N7gUQsReKJbWzgqf2ogGUqUQs+5JO6xr+cd4rHBnCyUga9ktuN9b2c4obYFJooGSeF/RAKhb3p26eVeiLwLjUJMj8hHmPQZdemyPYpMZC9xJzKsPBniQd38BihPa+q60jLNS5FhfiFX2lQup9xe27M9KngNYsTfPlGyCGa9ERA/uecLBBR/y+oj9lef8D9XK+gQMvUapiLaRTysUJM6cf5CYcCiGmHINy91iRg9inBSEwdtXiV4gPFPpsH1zek4hFD6dONjI+9/xYR81V+SwkZgiHBshz1GwcTA95Qx7+7sRLx7SMMyt7po1fbj7NgUzHgYHfDq3mdL9hfVyKWG936XRq1p9JcyI3KFzZLbm1ipmPbjbJ0BwKqT9wscOnxxGU9JarDk39a+m/R6GY8ZYQATfsBW0llszzTAlUhq9/qVSIfDpUlwHLWn43Pw4B88UOaxqMmGhxwug3R3zsAMdFNVfbCYLI4sdEAna2SGVFBaNq+VFJQoT2NPZUSJD7RkmLukV9+ofTIJGK+leoLV+Nt+jFXWlFsPl931tIxAEQJWC20lXOF34xRk9mxv4Ihoyu7cflbNascdj1usQ21N2rRDd7579mN6TsZWP3tQCB3s/co7VpeEMb+3DIf4uxy+jzPrnlssZS5XPfmBpu6ky5h3NLlmqNYdQvUooy+Wt+5GJssRZ4WnkUGlz8livaWEm1Nz9RgCvoM2cp0qafxsYbVRuGlRF8GmGJW9KwZ0ENWziavCjW"
`endif
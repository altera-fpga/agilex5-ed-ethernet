//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vLW9upZF1KgEgGonSIM+HzyGLuor9ej/HbR6O+YHtYpBSJspQWExGFpSJYg/
krXV2T08qa0omiqbjrMHzerNcdilVNcwOdf3p75w/4WbqTMpWN434fQYbKdU
25tuhfqczwldA0os87QnG9XDNGyP6oajXsaQCfXUy32P14mBiybSNJo7iM/z
iwaBE/xslbI3e7ErOu1U92jc72Ymi2d9KTonLpNAdJV18g9uRMlwt4FvO230
a02Y7mYU+9udH07uhQ61dE8wjCvY0QG2fi3uLIML1H+gU+PJPqOdAHZ9vTAf
4xvZdzKHJaRRK8tNxjoo9YLFqFVvw5xQU6adxhPjkA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lxVmEM4Jc4j2HeZguJKnWpdwE6zMSNRFyV1I3eR/wqiYZ4Xloxa9blfvqRo6
fUAePuAStnUo9smHAviPQ7G2Z4DgTrYe7eCHndoMxUVQH9l9nvsTipn1DW1j
4qxe7BHwoaI3aRvZAVgR/jAiNTHbx2pqIk17nBpPhNTvPIEb9vZBT3dXibfW
SIrE8YNfAUENpHspaRGj97dq1CMYRQZAJuF2SyI6cM0BieLCd374kZ9Z9AJC
znQWK0B0eNQyfSjmA3Gqvi+FzJnn4CFH5858qeNZaTHVZvshNTmCmDHNsvcJ
FJxuh58uQ7BKVPadlqnHE7RVFFBhLk2ySz1xmuoKIQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BEFGw9YDjYUE9g4I5G+1vmg7KiAAfQNagDXHnARVwWu9NQt0zt18b7v/AscQ
Ye5nsEcGDyb29vZXb49AdzOf//o0LQGQzR1HanAJeB6zJAgRWca+rjH36LI3
/NNVUKp0wXptMjhoEYGt3uP8icmrkzcPyaCgz+u/Rgojg/asLHdq/W+8CQtD
U3L8jFkNtyuAmqZyUVkG6GfBGy1LDQqj+lj2xZS1h+7r91RtjIpHXL7OPjmT
0p5XFRzBWxKqWE7tvpkDSJJ1cD/fzQ4yHintqK9z3zMISNwZoX4qz7h6HA6J
bX7jg23i8w15WHWYpGZXWASlspe8T8q9OKFFpr2Tyw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YbofQ1h4YMJqfvr+eo9vryoW3+/taCF0D/sDOWADX6Ln2u7lItDkOaEAJAf+
AKdiypwxE+ucKLWjORQ2K23ZlsporQLNu3WEmkOmQwnbKvuZtVzPLXnr2RJD
XAgh/fVylxkSUpPd94MD6XzBFwc+X8rB/jskX3+F7jtvWX+sOsxP67wvzKR0
ZZCsCDua7CSTIk5Y/PnYXwb+P/wB3pBbAvPh6FoePdChKRCoJaozf2+A33bH
f1+Rq3Gc+dQ0lFGEQ96jBJ0YUtoopOwzqjIVkKTrdSlO/Ct7wVnYEFOV4K91
Thy3k+MXbrsA7b+unBmeYcH/AOklJopMSnfLxHzIvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OXHElMMFEuIFq14x3oHpxei+NvVkSOb55P8+wONkQdGsYNxV7u1WLfXTSO6m
sOIaiU3y4T6LxkOVDJ7UF0KA0SIQIdwOSM6uMvugTDPnDjs4xQjZLH1++Pn/
bl6TK4EwOe5iE1RLve5q81N5I8q+xe730kxXSSEB4T/7Yqa4pqk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PFh7FQrEFdDZtglS93oxriHFEMAUuP4VJjnI2CqRnm+/NWNjTaNVsrYeYlLc
skOgF/Qz5LtON2sUr5sUFRA+Q3bP6EUWkQX82O6bzp0u0BxXoQjKKvofO2vh
j2o0F/UqeTFkclDg2WvgbEfLbNOx4f2xtkRvSF+5BzyI0S+BbQrtGWqRcLFy
6usjfkLTEz2cVKRbha1dqkJvCBblS5cFd7DhVhY/ne8VIc/+JfLj1cDrJFWT
riZOFiZnQR7eHtGw5lIUVf3EZstHiTsD73fZBL41WsQM8AnsHG/e+rFzkCEQ
CKceolBF8CcJMljtl5TzP5Qlyf8PLJXMksjTe1LGQ1CopG7+CfFL4z8N6aS+
jpY8kHDBeI0WmGWz4RqQzMOavJl1odG85zWUn8B+NpY89U+BwQnhkrl08vyy
u0js1eIF+hCTyhqevJ2QpsC7lz/So08vnxZrUcKz3KcMpeKzi/0gzNTQnFEY
i3hzD+4ZSbBz4oW7q2vIqngdBI9kk690


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DtOiuJfCbT5QuRZvv7QTUFuPZt00gk9S63yXgQuDZr/eeY9ilbrZ2Bs/aWAB
tTwum6vsEbukeTYaeppNQYtMT48B4c27tmsB8ATHx2wOml8K4blfT29s9ULy
u+UPsHwk2TZturc4zcToeZAEpHsjXedqM35R9yFom6bRYi2KsF8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fxoYvJj+hHYnWGASxARpteEDt04VcufkpuPtWobdMu61Utnrb6AoVuekuuGq
bOtfCGFp5fe1BNVvb0DvjaljauEzyHaxmEEVkshjTEm6mZQdf8pgSRGB8PP4
6qRQwXP8D769dXgzMlAcGm2f60LobFXwDQq0xlXq4xhlYiYOktw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
znc4Wp3tK8iA+uxu+SBeqdSRUP7h1OMPYY9mzvHLzf/8lPDFXKa5WRLyT/pe
2wPSrlbwh/CEZoNwlMv9EdKJS6MjdqSCXpyCGEmhlef1cwUPj3EzfYUccOlE
VoslpP1yNLbDfM2yiEL7qWNd8OtJmA+/QGeSKrRhs9nbyTC3KNd7fJo149gx
hzOCvqVf02EdiRkxNt4pC2FOcXM2K3v28Z/Gtcc6W570eINIuOYGJK6giWb1
KEbJnOJWQUqgZMLh9RlG1m8WdEF3zAhx+gt3Oy6b7yf1LMHb6bPENMwr/3Oe
hLiYQe6pNS+k/44Yzie+4HIOCxkEnnbkzLDcN9N9eWHe9bPfppSrGRWQf8Gc
HMeE6hN3m2VEPBDQhe6odBgbtSWSOKIJwTy66Jgq4kH9x6Tz0/E2VTKZzBIv
y/wlMrJKqeHNPc4TswI3AHTKrGqPEb/wCdqEUdhrS5g9vZz6DHRYD+JRrykF
sa+FAMbmw2YZplDgFxo1zywXw4GKhvQQnPonoJWsKSUp2CQPt2yq2rsp0Kqu
5Wc4hQ3zivTeBjVlJX6MY/DYfTsn/fCFyPykZoTkXrEXCYLR/uKFeSF9g+ko
TkUJakPLJy7kNL4E6zhCR2AxBmrtLZ6HrgIx5TGBF00K1WKYF00k5//8Y+2h
mVWQcjrSAoxpIdynM9qCDr41AjXFcYoxfqIOoI3xWLeqDiBbGRmRR/dP3V4k
WgghyIwhB286OexPNQXBU0aMuxr7l4/YpkIQKWTUQuFX/tI93/vStFBmBbMT
DSASHJ0Hv2j9WguZ+n6iUEECu2HkJDmgwmqvR4IL+R06AtezcXPxSl5rlIzo
2oWeThe2XggDXlB1T4kEnlIwYNjodQXBguGD61K/j0EXSzzJpBhwKnb1/Y3p
9qPOrrRhmOg2Wuh+bUlTIVCFC/eE0resJhvcHw9nSL/VW0/u7UzoiSDqW6Sp
FlYys3y+opPhKSiVXmp98udgoYq3ZU8YKCK++pv6ofO4b9xpVBmhply9AKIU
jwRUuASg4y21evr1r2ub40G5iE8NsKvD4hIueXgy4v8x+EUcYEz1OetwDUq1
SHaqSs9LYsJTAMEzu8e1c0pbMA01h5yoQfMvXDD0lcYukBKhhF36z6jcOU77
EWyhN3P83FuuR6ZgESk/ET90KRFllNGyvN8mHPocpopS0FaM6S52TjoNNhEs
eU3Cvo1rn5Fs16wEE4y8VLesY2+hXDcp18qc8MA91AkLS8CXY51weEGYTww1
pI+I2rmA9CYSEpq8oMV6P2snDcSkfSCCmUi2ugUWLgcOL2Y2QdyHrETbmY5j
h0J3Etwy6WzFD1cF+eLfEOP0cmAo7LDUGOv3Knz3qBTx1rjYoYGTKJR3bUzr
6lnSi+FahIMS8FKIh9Xdlug/gYKJ4otpVKkiwb2oIjAlvsuY/9Dz8wHNB9GZ
e/Svj3fHtjsl+SNGoHuVgnh+rXVGg9Yvxs2Lw+xhJW65/CN0H+rFznAOyh6r
H91aNgPGJ4lxOv/RyjMyi9r2tQZafV4f1KMaDUDIIWuEJjzXljwrRvl4UYNG
R0fJ0TdjgDA2RdO5DWeYL4Oo+2x0s7qUPvQGPN5vPP1+ABKAdbOHKev/A1VC
HETLWZCrDhEFhqN1fSY2P7AMfHleJKu0kEl8TOxlvp4VpMIW6pCnT2v9cUr4
FiQfxtuLVAOv95Aoo29qyjKnYLZGlO7smOuFEit4X4lCw1hg+DwJ+MYTaDnf
0DZUMnshnoCUB4+CYi7GpVY3VOMCyCkA2tVgfcE/QInSXaDcHBcwtVqt6a6U
QOy/mE5ObZEUzw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI39S6hag5+m5Z/spi6cyCheh+iqP4+n6Tm5wqzlkWJLD4KnNyQ3NFg3UFlQte0JZgn7mHwJ2Ujisjg3jYhPJN4Nyn8F8g3zhaKlg1W5RTnr2zjcH1a7uilMdnXt77N88SeXlhjILebSc30RHmFcaqktCR/j2XIFSnfKmpzn2v62bQ/n9MwGXc+0CtT03E7oDHrX/8WPQS3J/WWSS90DBijapLRBEPP0MkkogkemPfnrNEm+iTa07An/NvYO6yZxx5HRvRkdcDiG66F2UGgBd63CUjGpiSxCb0u1FOyUVkeXG7yrv8HAYwJ+FMelmpqWz+hxuNYvc8o12h6BUMaKr4QEJumvwJK31I+6Ns0krOmJMrEG7WwhcRVHqwzGnCC0jTMNIJXu3aBi1bB0W9KqqNgOllf/zgH8t9BoTyorwaP+DkccJCqqrE/Jlj0DssY+8ct4BDlSyKINk8N/S1viA98Bat45yI1NLkgr4+lk09UHBpZRC2Mq7HLDGbV75b8kof/2ZAmfCypUEzTjfYWcHW8HZr97FzaJZ2Xvtr2yaUcIJCPjqIfxPzbJWrbB8pSBdG5SictWw3lWGUG8h8wSRgg/Xd2p0DIc6sE9yicFlL90Zsynlx5nKpBjXVZTcomq70k2xK4sTcW/6I7Q2TtyH6dPO4Hf4zTE4a9jIpuFSyN2LyrVXjbi/QtNOrGI9Wz+RlSjPY5O/wPHz48dC40MxHGoJS4PjTE1nFfofeQ2EqthNQKeN4HN8bWmp4cXW2NOUW/Pceqh3s9oUiaj1SKooC7z"
`endif
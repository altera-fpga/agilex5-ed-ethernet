//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bV9fDS8Aja5XSd0AJqhsoAHui7lrQmOL6SBIolPOBqRLuoeyPnmE9W03kp6R
gUiMAdzDYQuf/R934WpaThZBBXl9X+AdPZLrr/ejeAG8iWXMh+7xoiLZCjij
AjKbTfGGwIX3Duivdo7ARMTaT/k6Rt2xIIH/QDu64GzGhcLz9QwMW2p4v5Qi
raOx6mVbXiPyPKfPYr6hTVWnZ+IjkPLHWDotL+3D+MvSuMgubkxCtbImvIwm
2XqkRD5MLdoR0j2N26Hs8zQcx22qtiqarVkFg2yuZKaHqbmArVfAkETWP9TB
gcjcv/SQW7A6bmZGBGZ8Y2SxKeN0vc7l6bRuaiz+og==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ozBYJh71xdl65cEPDcmDj9zPArjfTCzOUL3eqqyvFD810hiCohOBwRvlK9Nm
sGHqs4LEkCHZMxRObaX0+aVqaJMIIGJOhjrgGN4H4rYMZXX7h86e6cpVWqyN
Hp5fgq9TK78N9LSYjzsctUCdE99b0eprpPs15xPSd1BIlz3i/+7FOKH57P6Q
nI1ufP3hanBqA89ext61OduMcG02/hB7jveWT6ctnpu+tGYQLnI7S3izP4XB
RPfW/bzFq8LMrK0q34Sc6BlCypPsa1LFZLSsxSBaqdFUVydNEh6iIEtLlExC
UuAUU4JKW+vzx1wjuQRpRH/hjjFe+S2BNFuXcBdHQg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b6Y/xxk8yXVUxu/s77gGt1aVyJzji0OohL1DjP2ETwMwafN6f61rZOnZdFCp
WE4oEqZeGuM4zgBaZ/5G+JdR0Lm9ubLMXCM7aqfCCQZPBeJ2VqLIFRC52/Av
f6gZIxK/uW47RDi7jVpzjgqyCF53lunjWyhpdYNCPywl32k/aWCeNj4VOI2w
dKEk+U/rfT8e3EZUWCzPL+dV/VkMjeo0TF98uHZVofGApvZu9izch2Z5Bvso
ZKoceyl0M9W2K7HcQxOkooALhp7aDSOo1qe5ZXhXpDFmfzIXej9XJtOY8cUU
VFqu77YaA7uDVxojWPasFAsA0kVN1DadMXHg/tCpJw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hikuV9hTYdIkXXmyqA+BYyiWl+LVgHXqQq1mw74jwv+YsW3TwIp/+liMGLxd
HiZX80bfXFxiOnfJzYb+gpnttNBObcY/K2ymkYKPiJ1jBt9WExlVk+BjIHeA
hXKaX7bb2hN8ASywmweOzMPxhzDGDc/pXwE7p6BQxnc/Sn1AGvozQcbx1vtd
VvOfRRd6jPyHxa0rd/X7fZOI88QaWtRv6tij4QbF15DJqgcSNrfAyVl6ORPw
HdeyJbc81QdUgsXqiCdqvb6qUHk5Ib8DWDZUnk7sLYSWkpXIzMcDRj5GgK2j
zwgBovD5xCBalFoG8nJgmiBymBOjvX7wLcpYtV/rVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r/ALBs0wCsbcG8gmyFGBkd73/ph3WRw82J+YOWzitPd39nlsLLYSHLFxL3j7
nzUS8+1SZPY9TjDqu36kvY6fIiNaKMkyJZkTiXgBq32o3X7gZ7OH6NRvE84i
EW8jFteTSdXNGMZu4CehRJ8GnTBRl79/88OUOomFZE6L7XlLjUY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HNchphLwALlHsM3ZOGtN1cHL/xUAIG/DkvEaPKtzzwoRmDMEbBNWHFfEFdx0
GuaF+4WCZQsRe5oTCuNUZ3LkpzZk44M1KJuAJr8ObsMCckjKI6+kOKzU4M1d
7dsgOaIqrda2kiGIwme0uT4aApyI4ElU5hJHIeuxU5caOB5Yi8uLadvRoaCf
T+R1foMLE65vpdLZ5TWQO3MKw7eAappm3cjI2rfQOVAPoVLaGK4aVe9hGaRU
2T6/xmi+1jSN0o6HfdqxNGSxkOBDoGT9Ngh0kfay1g6+l60b9YR9HCMc84hX
0/2YQsik8MSRdccdww2fITgzgGWBZpu/vVwD4sHNC84RrlnFMrlfDZGdzP/H
W4RHv0EpEh3cq1is/ao8rVXRUDglOAtth1GiiT+Fug+tpbaZDBlLo1rgCTtR
75/tiylyT6nsQz2UA0fWKPx9zyzUIhvXx07HPqrdt0MJyBFr3tGiuE7rFNzS
VCq+/FWWo+2Conqhfu3pr8Tf4w0zGz6h


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z6nk0A9GaMWJF/MzNTr6ehFlK50yXKSQlxYldr+SbHuuJhsroXyGPpzYRZmK
KzTjoFUmIxlphPZ4YZqZbRMKxZ8hGFPUaU97Xk8C4FztdCcqVPLXxkn9REyA
rckqVXql6LglpL1y7ve7EvMCCZe72l+I9CYCOk52MaKrwjaf9iM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iZdMElQ4PuPRzV8Yz4N87p8b1mBLEXJ8HrOEPzu0Bb8SSe9JBEBWtPdwDX64
pFkUnEzzVhUoKQ5LFt89waK3APL/ed46Wg+U+RsKITkCFW7ToI4S3sUD7yWA
4m/iJ/6UB6MoX9HzrkyR/XSKtj7X6qT014rB/LC3cPLfTm6jRBA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1232)
`pragma protect data_block
nL/XWe5y2RVSG4OeMHUZRIagoJN8TP6tE65y7Gd2rqClDlfKvGHAeoaAApyj
15iRvYRKwwELRpRBjR9Eox4+f8nkLvu34/ahQsaKiK1/uvLB128055vZEYim
jU8/x7aerI98aN1vt4LAJrzc30b/Rg/X2XElqKLoEKUKibrEFEQPs89NqVp3
mVzdpAtVseHQ6WdIa9jsYs0m8iss95YJbAU/53VKo5XS52x0sJc378i3/mCW
xyLtGkRx5Udc8Oa6J7RmGNl0Fkvb+2tvdIxxRNHaTKCSt/InmfRe4rVJdz4p
q1AcG7KBRPXNONEQFFqEFlvpBoik1bOtRXiL/qjPKoO3w7839NOu7H9DcuB5
pPo54ErIo/9oEpzfmyfMQJ50YL3ctv6+U93Ui4WNHO6xKi51esw0R6pCW0NR
EJeszS+1+UaJZjd6t+HRl1kFHqtV394Z9nsb/AoQl2XMsqkHGAoE5l0O5hSb
b/mOI1zf4hUJiP5O2TQK30pzxyxOH5RL3e5B2phOJUS7cKcp+S7u+I0+aaaY
wgfOpvt4ulRJpYz8ZfBVUDNJw3Lzp/m1XUkHdctZp17oYhq7jH9/iVOdjieB
9WxFKDnvp+udNUFWy00Y8wTzzVTKHw+HrlGnsAoyadvSEdhdrMco8qf2c90+
2zHWXbYoXCVV8XQQfZE9no9GjeEWUhFEV4WokVKLaOfEgmWQpm3TfZlu403k
qNBVCIJtftRkHIHaLt3/Dc1v3/WsPW3PT1yn83jBNiMmjKDIR6TJaxEtmAXr
jQt9VxQcdPt/08l4HcQVIKjofkAzyJ+A7Zyh2aCOXUvWDR/yW6JqyJGg8PDd
vGzIT9FwUqzdidRUmHRUY8U9aAnIxDwbBHMi6TtxgCpmagjDsapF2z3Vtubc
8xYGXpovmCFSI6DgXPYaL0RFlEJlA6lYkvXm2J5w5XasNLrM5wzaMNAKJu7d
Cg1moQpXePG9vPUc1whowXyWfSu2aVw0JU8OpuqJ4EcqFoc1z9rjP8uyUGm3
Z3XQ9swqxRBB/mpNXUfKIy8sm271KL79EPWgeq07ro/cC8GzsBbEKBVuJsIq
+3x+vrBbekRtLj+KNqMsl+6r1Sh+JJypYp/c5+H8K95fa2JQCmTGg1pLohon
5m9jwLcZdzkIZ8DbBoECe217+Yk7RoZPBV8ohkMNOwDG1dtcDX0ZO1fOmtDa
YCfEN1G/rd/iUBSiTxGRzypzqy0ZcI0Fj2YppI9Dw6GOIlUAzaexDDicF50w
q+9XhBzwJH0sycbvy1jVIquRUR6GhNF8nHLKj0b/6r7ueJ9G+v/y2WQcl9Bp
r0gJBWkoS65+8i58ffIZZQtDWeVK2L2xgXbg6btyd/5p+J2/UruBcDfEp22a
1YqipZOuMf+uzK/jRKgjw3iKWdGuLubyX/N2F6ogZVXMS8kFapNIN6rG8KAH
ah6qbWKyKGUvZPLcg0U/WxwBS5pGKCx/Arnn6XmL7tpIEzIO9wtjkWwjDEEs
24tXabBqUa8s2YEld+UUKjbhb4hASl1uCjeJAVI8BXimu1COL5MYF6hvIiKs
IsU048SOXAKNTMIvZhpnhmLp1V80JCcRkJ9QjjIYlysaYKMRhUa4f19ILcwp
fXt9bWs0CnW2Oc/y/iTsqZU=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NdOh/z3LGtaoyYmSC+C5BVVnr0UAb1ltTHwAhIFCaqEz6kGoYkY6ediorH+Pkty4P5IckEz08IGB28/SMfP9I/PHMhE9lbJVYr6R4FPCLMzhT91Lo735SBGekk4rkgoebNeUyj8aY48r+doq6izRITr0ceVBf5y4K5Q93CbDlDhY9IWU8HWRKms01EECvSlyhl5r6DrDKQpIJvLOC1oCW6Iw5ooE0PgmnqlRjlCA/er4sIr+LdiaCAPrhyhrmZ0rgxbipnYJ6pX9ezPOW2DaWaOcmq/TYcOeYPLa9iLotfwyMp57h8x6XYgf/M7eeji5P1V/b6bqlI7tDXebe37InJzsFXTsaCruY0EXqO1H384u3Rbmh8l0jSpY2EUoZ0OiIwt5GA87IdA+2wXnTBC4etGTc+QW1VHDvW3iW/cHs3T5n40on0gOhPmTKECymWatzhWWgKgVkb+ugL2qcp8T6s7AKtUuWkOeV6qRpOgkZF6cP9WDV6oULF94n949pHjKOOmDhMwVTgbLve1pOXRajbntHpLb+J2YoblG4H3tGpfijz36tgvT2pXBjBHYxfCf7kgw94XvsaWqhpWtAEnnZZ/dNhXGJIeM9uM5LNow06i7t6LzMQ7m5Gt5hlR5XsGe6lWJiagkAwXyMKD5RPPiSTobfFnB2vqFdkWJYdbfvHuR6gyJLmo+JS/utR8hZSAYLqJI4Za8nduuGu5AIyEUcdebaqwvAMIA7fS8nyXxTsWdvk7ghM15GOpFETWxM72E+x3kI52TkMFgY8MhTuA/YZSVM5e8Thz+n3hxzsmuuepP5bnkl3pO7EhWe7PeK/7rl4IBnWRFjLMq/TMEFWTxVDj/IPmsumDY0DlMUcEo6w8Pic294G29bMkwaA3JYH9Qgodv++Xz9VyJ9ArItObpqGzxWWQyJbNem3Ae8YiARCvT+OQ3pjnotO5wHBPJpo6ZytyDm+IzEFbT/m6WD1+gkmKOzRsxO7OBQJL/s6uvYe7riubkFhJRmUY9miTqY1/G"
`endif
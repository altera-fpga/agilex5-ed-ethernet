// tcam.v

// Generated using ACDS version 25.1 129

`timescale 1 ps / 1 ps
module tcam (
		input  wire         app_ss_st_aclk,                    //       axi_st_aclk.clk
		input  wire         app_ss_st_areset_n,                //   axi_st_areset_n.reset_n
		input  wire         app_ss_lite_aclk,                  //     axi_lite_aclk.clk
		input  wire         app_ss_lite_areset_n,              // axi_lite_areset_n.reset_n
		output wire         ss_app_rst_rdy,                    //    graceful_reset.rst_rdy,      Graceful reset ready signal from CAM
		output wire         ss_app_cold_rst_ack_n,             //                  .cold_ack_n,   Graceful cold reset active low acknowledge from CAM
		output wire         ss_app_warm_rst_ack_n,             //                  .warm_ack_n,   Graceful warm reset active low acknowledge from CAM
		input  wire         app_ss_cold_rst_n,                 //                  .cold_n,       Graceful cold active low reset to CAM
		input  wire         app_ss_warm_rst_n,                 //                  .warm_n,       Graceful warm active low reset to CAM
		input  wire         app_ss_rst_req,                    //                  .rst_req,      Graceful reset active low reset to CAM
		input  wire         app_ss_st_req_tvalid,              //        axi_st_req.tvalid,       AXI-Stream request valid
		output wire         ss_app_st_req_tready,              //                  .tready,       AXI-Stream request ready
		input  wire [7:0]   app_ss_st_req_tid,                 //                  .tid,          AXI-Stream request tid
		input  wire [491:0] app_ss_st_req_tuser_key,           //  axi_st_req_tuser.key,          AXI-Stream request key
		input  wire [18:0]  app_ss_st_req_tuser_ppmetadata,    //                  .ppmetadata,   AXI-request packet processing metadata
		input  wire [0:0]   app_ss_st_req_tuser_usermetadata,  //                  .usermetadata, AXI-Stream request user metadata
		output wire         ss_app_st_resp_tvalid,             //       axi_st_resp.tvalid,       AXI-Stream response valid
		input  wire         app_ss_st_resp_tready,             //                  .tready,       AXI-Stream response ready
		output wire [7:0]   ss_app_st_resp_tid,                //                  .tid,          AXI-Stream response tid
		output wire [491:0] ss_app_st_resp_tuser_key,          // axi_st_resp_tuser.key,          AXI-Stream response key
		output wire [31:0]  ss_app_st_resp_tuser_result,       //                  .result,       AXI-Stream response result
		output wire         ss_app_st_resp_tuser_found,        //                  .found,        AXI-Stream response found
		output wire [5:0]   ss_app_st_resp_tuser_entry,        //                  .entry,        AXI-Stream response entry
		output wire [18:0]  ss_app_st_resp_tuser_ppmetadata,   //                  .ppmetadata,   AXI-Stream response packet processing metadata
		output wire [0:0]   ss_app_st_resp_tuser_usermetadata, //                  .usermetadata, AXI-Stream response user metadata
		output wire         ss_app_lite_awready,               //          axi_lite.awready
		input  wire         app_ss_lite_awvalid,               //                  .awvalid
		input  wire [31:0]  app_ss_lite_awaddr,                //                  .awaddr
		input  wire [2:0]   app_ss_lite_awprot,                //                  .awprot
		output wire         ss_app_lite_arready,               //                  .arready
		input  wire         app_ss_lite_arvalid,               //                  .arvalid
		input  wire [31:0]  app_ss_lite_araddr,                //                  .araddr
		input  wire [2:0]   app_ss_lite_arprot,                //                  .arprot
		output wire         ss_app_lite_wready,                //                  .wready
		input  wire         app_ss_lite_wvalid,                //                  .wvalid
		input  wire [31:0]  app_ss_lite_wdata,                 //                  .wdata
		input  wire [3:0]   app_ss_lite_wstrb,                 //                  .wstrb
		input  wire         app_ss_lite_bready,                //                  .bready
		output wire         ss_app_lite_bvalid,                //                  .bvalid
		output wire [1:0]   ss_app_lite_bresp,                 //                  .bresp
		input  wire         app_ss_lite_rready,                //                  .rready
		output wire         ss_app_lite_rvalid,                //                  .rvalid
		output wire [1:0]   ss_app_lite_rresp,                 //                  .rresp
		output wire [31:0]  ss_app_lite_rdata                  //                  .rdata
	);

	mem_ss_cam_top #(
		.CAM_ALGO                    ("TCAM"),
		.KEY_WIDTH                   (492),
		.RESULT_WIDTH                (32),
		.PPMETADATA_WIDTH            (19),
		.USERMETADATA_WIDTH          (1),
		.TID_WIDTH                   (8),
		.NUM_ENTRIES                 (64),
		.BCAM_MAX_INSERT_ITERATIONS  (20),
		.BCAM_TABLE_CRC_POLY_SEED1   (389490449),
		.BCAM_TABLE_CRC_POLY_SEED2   (655828753),
		.BCAM_TABLE_CRC_POLY_SEED3   (757182871),
		.BCAM_GLOBAL_KEY_MASK        (512'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111),
		.TCAM_CORE_TABLES            (1),
		.TCAM_ENTRY_SLICE_WIDTH      (40),
		.TCAM_KEY_SLICE_WIDTH        (8),
		.TCAM_PIPE_CTRL              (19),
		.TCAM_GEN_PRIO_RESP          (1),
		.TCAM_USE_ECC                (0),
		.MBL_MEMORY_CONFIG           ("SHARED"),
		.MBL_LOGICAL_TABLES          (1),
		.MBL_OC_BINS_PER_ROW         (0),
		.MBL_OCB_TABLE_ENTRIES       (0),
		.MBL_BINS_PER_ROW            (8),
		.MBL_LOG2_ROWS_HASH_TABLE    (20),
		.MBL_ROW_HASH_POLY           (1637095),
		.MBL_LOG2_ENTRIES_KEY_TABLE  (20),
		.MBL_START_POINTER           (0),
		.MBL_SIG_WIDTH               (8),
		.MBL_SIG_HASH_POOL_SIZE      (8),
		.MBL_HASH_CHECKSUM_SIZE      (8),
		.MBL_KEY_CHECKSUM_SIZE       (16),
		.MBL_HASH_CYCLE_MAX_BITS     (32),
		.MBL_MH_CHECK_KEY            (1),
		.MBL_HT_RMW_EN               (0),
		.MBL_KT_RMW_EN               (0),
		.MBL_LOG2_TABLES             (0),
		.MBL_TAB_WIDTH               (1),
		.MBL_LOG2_SIG_HASH_POOL_SIZE (3),
		.AXI_MM_DATA_WIDTH           (256),
		.AXI_MM_USER_WIDTH           (1),
		.AXI_MM_ADDR_WIDTH           (32),
		.TVALID_PSTAGES              (0),
		.TREADY_PSTAGES              (0),
		.TREADYLATENCY               (0),
		.AWVALID_PSTAGES             (0),
		.AWREADY_PSTAGES             (0),
		.AWREADYLATENCY              (0),
		.WVALID_PSTAGES              (0),
		.WREADY_PSTAGES              (0),
		.WREADYLATENCY               (0),
		.ARVALID_PSTAGES             (0),
		.ARREADY_PSTAGES             (0),
		.ARREADYLATENCY              (0),
		.LITE_DATA_WIDTH             (32)
	) mem_ss_cam_0 (
		.app_ss_st_aclk                    (app_ss_st_aclk),                                                                                                                                                                                                                                                        //   input,    width = 1,       axi_st_aclk.clk
		.app_ss_st_areset_n                (app_ss_st_areset_n),                                                                                                                                                                                                                                                    //   input,    width = 1,   axi_st_areset_n.reset_n
		.app_ss_lite_aclk                  (app_ss_lite_aclk),                                                                                                                                                                                                                                                      //   input,    width = 1,     axi_lite_aclk.clk
		.app_ss_lite_areset_n              (app_ss_lite_areset_n),                                                                                                                                                                                                                                                  //   input,    width = 1, axi_lite_areset_n.reset_n
		.ss_app_rst_rdy                    (ss_app_rst_rdy),                                                                                                                                                                                                                                                        //  output,    width = 1,    graceful_reset.rst_rdy
		.ss_app_cold_rst_ack_n             (ss_app_cold_rst_ack_n),                                                                                                                                                                                                                                                 //  output,    width = 1,                  .cold_ack_n
		.ss_app_warm_rst_ack_n             (ss_app_warm_rst_ack_n),                                                                                                                                                                                                                                                 //  output,    width = 1,                  .warm_ack_n
		.app_ss_cold_rst_n                 (app_ss_cold_rst_n),                                                                                                                                                                                                                                                     //   input,    width = 1,                  .cold_n
		.app_ss_warm_rst_n                 (app_ss_warm_rst_n),                                                                                                                                                                                                                                                     //   input,    width = 1,                  .warm_n
		.app_ss_rst_req                    (app_ss_rst_req),                                                                                                                                                                                                                                                        //   input,    width = 1,                  .rst_req
		.app_ss_st_req_tvalid              (app_ss_st_req_tvalid),                                                                                                                                                                                                                                                  //   input,    width = 1,        axi_st_req.tvalid
		.ss_app_st_req_tready              (ss_app_st_req_tready),                                                                                                                                                                                                                                                  //  output,    width = 1,                  .tready
		.app_ss_st_req_tid                 (app_ss_st_req_tid),                                                                                                                                                                                                                                                     //   input,    width = 8,                  .tid
		.app_ss_st_req_tuser_key           (app_ss_st_req_tuser_key),                                                                                                                                                                                                                                               //   input,  width = 492,  axi_st_req_tuser.key
		.app_ss_st_req_tuser_ppmetadata    (app_ss_st_req_tuser_ppmetadata),                                                                                                                                                                                                                                        //   input,   width = 19,                  .ppmetadata
		.app_ss_st_req_tuser_usermetadata  (app_ss_st_req_tuser_usermetadata),                                                                                                                                                                                                                                      //   input,    width = 1,                  .usermetadata
		.ss_app_st_resp_tvalid             (ss_app_st_resp_tvalid),                                                                                                                                                                                                                                                 //  output,    width = 1,       axi_st_resp.tvalid
		.app_ss_st_resp_tready             (app_ss_st_resp_tready),                                                                                                                                                                                                                                                 //   input,    width = 1,                  .tready
		.ss_app_st_resp_tid                (ss_app_st_resp_tid),                                                                                                                                                                                                                                                    //  output,    width = 8,                  .tid
		.ss_app_st_resp_tuser_key          (ss_app_st_resp_tuser_key),                                                                                                                                                                                                                                              //  output,  width = 492, axi_st_resp_tuser.key
		.ss_app_st_resp_tuser_result       (ss_app_st_resp_tuser_result),                                                                                                                                                                                                                                           //  output,   width = 32,                  .result
		.ss_app_st_resp_tuser_found        (ss_app_st_resp_tuser_found),                                                                                                                                                                                                                                            //  output,    width = 1,                  .found
		.ss_app_st_resp_tuser_entry        (ss_app_st_resp_tuser_entry),                                                                                                                                                                                                                                            //  output,    width = 6,                  .entry
		.ss_app_st_resp_tuser_ppmetadata   (ss_app_st_resp_tuser_ppmetadata),                                                                                                                                                                                                                                       //  output,   width = 19,                  .ppmetadata
		.ss_app_st_resp_tuser_usermetadata (ss_app_st_resp_tuser_usermetadata),                                                                                                                                                                                                                                     //  output,    width = 1,                  .usermetadata
		.ss_app_lite_awready               (ss_app_lite_awready),                                                                                                                                                                                                                                                   //  output,    width = 1,          axi_lite.awready
		.app_ss_lite_awvalid               (app_ss_lite_awvalid),                                                                                                                                                                                                                                                   //   input,    width = 1,                  .awvalid
		.app_ss_lite_awaddr                (app_ss_lite_awaddr),                                                                                                                                                                                                                                                    //   input,   width = 32,                  .awaddr
		.app_ss_lite_awprot                (app_ss_lite_awprot),                                                                                                                                                                                                                                                    //   input,    width = 3,                  .awprot
		.ss_app_lite_arready               (ss_app_lite_arready),                                                                                                                                                                                                                                                   //  output,    width = 1,                  .arready
		.app_ss_lite_arvalid               (app_ss_lite_arvalid),                                                                                                                                                                                                                                                   //   input,    width = 1,                  .arvalid
		.app_ss_lite_araddr                (app_ss_lite_araddr),                                                                                                                                                                                                                                                    //   input,   width = 32,                  .araddr
		.app_ss_lite_arprot                (app_ss_lite_arprot),                                                                                                                                                                                                                                                    //   input,    width = 3,                  .arprot
		.ss_app_lite_wready                (ss_app_lite_wready),                                                                                                                                                                                                                                                    //  output,    width = 1,                  .wready
		.app_ss_lite_wvalid                (app_ss_lite_wvalid),                                                                                                                                                                                                                                                    //   input,    width = 1,                  .wvalid
		.app_ss_lite_wdata                 (app_ss_lite_wdata),                                                                                                                                                                                                                                                     //   input,   width = 32,                  .wdata
		.app_ss_lite_wstrb                 (app_ss_lite_wstrb),                                                                                                                                                                                                                                                     //   input,    width = 4,                  .wstrb
		.app_ss_lite_bready                (app_ss_lite_bready),                                                                                                                                                                                                                                                    //   input,    width = 1,                  .bready
		.ss_app_lite_bvalid                (ss_app_lite_bvalid),                                                                                                                                                                                                                                                    //  output,    width = 1,                  .bvalid
		.ss_app_lite_bresp                 (ss_app_lite_bresp),                                                                                                                                                                                                                                                     //  output,    width = 2,                  .bresp
		.app_ss_lite_rready                (app_ss_lite_rready),                                                                                                                                                                                                                                                    //   input,    width = 1,                  .rready
		.ss_app_lite_rvalid                (ss_app_lite_rvalid),                                                                                                                                                                                                                                                    //  output,    width = 1,                  .rvalid
		.ss_app_lite_rresp                 (ss_app_lite_rresp),                                                                                                                                                                                                                                                     //  output,    width = 2,                  .rresp
		.ss_app_lite_rdata                 (ss_app_lite_rdata),                                                                                                                                                                                                                                                     //  output,   width = 32,                  .rdata
		.app_ss_st_req_tuser_tab           (1'b1),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.ss_app_st_resp_tuser_match_array  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ss_app_st_resp_tuser_tab          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ss_app_st_resp_tuser_ptr          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awqos                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arqos                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_clk                           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_reset_n                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awready                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_awvalid                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awid                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awaddr                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awlen                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awsize                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awburst                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awlock                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awcache                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awprot                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_awuser                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arready                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_arvalid                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arid                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_araddr                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arlen                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arsize                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arburst                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arlock                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arcache                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_arprot                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_aruser                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_wready                        (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_wvalid                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_wdata                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_wuser                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_wstrb                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_wlast                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_bready                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_bvalid                        (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_bid                           (9'b000000000),                                                                                                                                                                                                                                                          // (terminated),                                 
		.axi_bresp                         (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.axi_buser                         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_rready                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.axi_rvalid                        (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_rid                           (9'b000000000),                                                                                                                                                                                                                                                          // (terminated),                                 
		.axi_rresp                         (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.axi_rdata                         (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                 
		.axi_ruser                         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.axi_rlast                         (1'b0)                                                                                                                                                                                                                                                                   // (terminated),                                 
	);

endmodule

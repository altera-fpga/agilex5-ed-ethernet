//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FAPjmMqFzGsH6c1EDznsW6sEPdkhdXtP9y9sdaqKP/98GnRvi9Gh1YeN8yR8
2sdvItUT6fVGzgD3I6FjiZDDQvHAJO6/JPIh7Aj0cPzcGBXu/vRW3vEQj/cK
/wIn9oK7PTYpZKHifxHjhHWjiQWJM0c5TIvPtz33MnCsVU6gX5GRah/FaOVF
DaZj9DjXc8uwJFwA610IQ2u5Z/cH4ROSeQTY53moXEwh9WarqT3zeREhT6Rw
EevZnuX3DpMF06ZUT7ouOjY6dZHt/mtp7cDR3BbDV8hCtF90PX/NB0Hf1mmv
vzXjiSy5NkfB1s3M+sbsfNosDeNaLZrie9vTA7O+2Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A/do/Fy1csDcO50KERDkQRxgG1JjY0a3uH/ZupwwOYO+PxalMTeKUp0drDNm
IVjK82gFTKEr3nmWE+ANvkfOLWAFZ5LBZCSEH+bTEJIDxDchxIVajE1hImWZ
HiVCmiUifYQ4dlN3N44wEgJhKUSWRP2gEjc434OidF6kj9W4i263A2VTCSJu
nPX9giXAQojmqfw0kI4XVtQmtzDw/dlCOjzDkMJDroESXyAW8PamIPzSjxHF
5iZwfcCiBojbW0WhXHHZXS6nzKNBJbjHEUsCCiKxRXCZsNHRhCyrVoZSFZZw
nKN3QFGpytTBTp5Ui/Jlt3F8TIdnSVfnkLr36hY4GA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LnptZTsvu7PV7Q7mt5fXg6dLdQoFOfLs2vED3yAZdOMn4QEgGy9MLF07M/qd
HvAq//cvvNf5hGPoNO0levlZQT/NKFjCOIEWBh22u+1OeZxy966xjMMDOrnq
5wz2DPV8dIc5TXV6AE0PGa1uFGypYbdxl6DVzC0RcZCz5UzxkG4YbWJNBYix
B/jAbhCj+JbJKzc5VDYbd61zrVcR09x6IiL5ZyHS1NeGS1IKOg4oRLxNwFIV
us5wijHITr5foa7AcjNZG2j8kuj/9/9EJ1c8qHfe9vT2SGR66QRqUuOagFV0
xqxOsnA3YQ2wzM8bDfsxtZ4QGusVH0+52im125Og6w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VxsUC3lp+udjUlIUjayUtK2juFU0YDXPX+lIXPXmcSbnBgUbQpm2o3HkRVMY
17QInVikYXvkDEphpH8Nb7nWxVf2q5zrxhzWvGLfcHA4C53pN+4nChkx854m
XTwI8RAKkH4vcRO7JAXQNEF/jxLDC7fwMeLLwjJfZeXHrWURNbyNN8RVbed7
J9gjZvRz9t0sSSLds9O7cfrh1uAQ0eFctHO6C7cQzFBCQsKcDaRE41qdOEbq
q5YVUwuusaL0FH0k27lB7ZDU5lJ3cogbRrfLDE9SWsD8inWjvC4j7gHz31XY
kDRKixsXVxpg+hq8OV+s0CvuPdpjym0Ugk/v7UdXjw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YaOsQZkFnarWqf7V79gBQ3gQsS3NtkoNpsLs3ug1nb5MvA1i0Ocf+8Fgrxxm
OtwxIvdaGvslTyYxFAUCjqrH72hXYTAqR/W/cvl0CbIlC0bHM0Y4LbN/Ly0/
WRgfIlmS2xl1ZNKHqm2KoNfQoQsU1CxA8KOckBoyfA6PkxQl5Tk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UdS7LB1ilowflWTrF9FH+JGTuf2USabQBLTu7ePSkQV+d3LU8TaXMx7RIdUt
rAd7TkI0591QBKa8VFM+levf+L0o1uVd2WgvruTiRZAOWfEs6zwpY4GGRv5s
qPnCIw2AfARB+lsIGLqKABfvpomgb4E7UtSQjRLoTopLkbYqzaIKAYoaCUDz
RAaGReGqkh2N7srCj0KlBGVhCTvumKdt5jPWn5oPf0u6PwpLp/oa1+b70LHx
ITVXuqAD74cQI7aZ2VBshq3hM5sOoycNtkqeVGDXxBXhe/zHVhmazeTwtdpp
abfy9SgINtVio00HYZmQqm3K1LHE1rUIV42FCh5aou5Aah6/gfOaUK1xXG8b
y4XXFpHr/MV9xLC1l6Tr62YXcHv5cpakujcc/dE4MPzbJabC9eWwTtaihr2t
Lz2KyRpu+17hEtSyuV3/EBIQRve6AfQzKHrnq1B1IIKhbtE9wvZM84BtukO5
sHVF5eXfJWh/Kh+yInLOpfTSaJVKy1wC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VpISJ+MGXaS7s5sOAcLa3FCcchRwLeoaNAUuEkf5tMVOCCCn4TCaXkL2+H0+
96yRy1467U4C/Q6sOeO6UEqQzE5AehtvZR2BJTXYAnBSsgbOEvyUJm8RTj9Q
XMQp6mgXMS4/cZDmjZKOveOrkpCjqZzLd60nMVNToewTWQDAE4Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S6k9mZraj4aMkrZqcIpc8xOZQ64Qq+ns0mrXkZJyVe8CrSUG5FmoTmmd6jR0
pWkwFZ22BY5Uq+9qxzBwFGZrV/6PzdyFfgzCp7pA09aY8nekecIZqEnAiz5g
OLpJoN84pphhD1FSHXbKzh8qr2hiZdxLEY9I99j/qdeD41CFTAc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4368)
`pragma protect data_block
QPtvlVaDjDnjq2Ur2Aq/PMen6satNKNtDSLuIWNxxjg0hzg/TFZb+BFSnu5R
cNKZL0kD6PITLMGLU38i8vDAbvzP3ic1xpIGuUHX371y9Y9Gjwqs0TWSueFP
oybIjW6qdmCsSzYKGIzEWiQZe1Xa14N/B70VfKhi6vD/rZa39VknYC86Ghuu
rheQFqJbZsypz8cns0vXVgU1bn9vPt6HssZhy4e6HPAGaU7RhOXYFREAWS61
xKcxvKbc08Csd298LaXgejCoyrkc4zWA/g+Tikvz73RBUw0M9ii9PuaVL4tc
0cUvWH4MCIsOFYH0+JBiAEACLGNz26psgAzQRSoS0zY/glig+339lp0CmZAs
Qu5gUvQrvQ60e7vTgx+19SADsQF2jhbpBpMZ7cQzDLJiM5MCWFd3ZjY3c8eM
+0z9QDZp7rQK/vPy79nL1HhZEyC31f4C/WI+lw+CSLFQ84Rt+yOxEqh7QPhJ
KEAbAcQDwBaIkiP1VYlP1KEc2vkRRiQJHN6F2cri89QzsBHo5I2UIYli0aF+
DEaKDXfax/weX35Aun+yqo1yH4tZAT6VRFjntp5KkkKZc42FeYYg/9QDypo5
9hqvGjsXhjNsI4LNUFF59Mvl3X6U+9Rgn0BVd0Vy0B3iJ0W5pd/D9tf0Byrg
J1zTHuXdd0+O8Kvh5R46jv+rTJ+iXAUt0GxsGfuVeYpqDx81Uagcbq9e9YSC
hqkDrquZKfcyl+HKzNtKtNPF/BPFZ6meFh1NeddeKV5fNwDcK9a3V/6k52NY
CDCNUFon4iW656P/TfYG9iRHokwITsmIEiWI3LR2xYSlUOYoRqBKDrjYhcLV
ZJPgaKGcQJ9+Ln9VE0xhVsaj7w634RmGKxXToQFheEmv2Z3/xS/iRuDyRSJ6
qhf78TZ0D0hUzFD5uYihF7sCWkb6O08oip9z0ISvyWQKrawRfFfUGpqqpqwB
3gXOoH7EwVaui/ErOxOn8cIIuMvrcx3/45HMG2+1C49IQ3IXei8uB1xHM9bi
QpKd6nDeBtYpVpI+4X90Vji5lBWyIwa5ZpsG8PncAE7suLiMzd0D6MIKLNGu
AhvqZrQ4BeNtmgNCD+31pIf8IMRN4usxe0mA97OsRielkgQ95XerI7Y0teMQ
R2Ub4xySjkkcO7D3UBGL/m6A/cPYCeRAYjnbVRKci5a6PqnFAF3bw1mPpmL/
820J4XhJcXDfL2f61YTFLNKXZG+ABc9P7b4PI2BYohTIfBKr7JDfUNI85tD6
Ll1IlVcFBgLB8fUq4nZJF68I2hhn9iDAv3tPXQgVJMZoxoCInTyNlWHsaBBy
l/Qyvh3fC9JQbtISeOoIs6MDQrIz+Dt+dF1qZ5DFyGAEIHgUOEFk8ej/hjxU
Ti0FpUdxik3btn3f5IdDg4gECqAZzMiNcRXrBFK0GIu90tBapvsnwi5Zb0Mz
lOYNCbC4ug50E1ONzabieQVn/yL0b+L/1lH76YXsZXx4e0S5NmbpChF6RGGv
ne8tfYR1mRTXOXZApkFYioq7N7sfFr6Q6G/DCoCxAeeRaDF2FlhZPpeEiaI0
w7Hq7d3Vy3SEBUk216XUaokFI8aEuThyvFjL/rzlVmxzpUerX/LF5bHaKOs5
oDU7+YFcQIpgWoVrD1RiRU1bnNahShjbdAgEZKv4Kx3bRyxbvo173+GRx9vO
9HU+6YxMTKqx+BhdAxCH7D1yAk+JNmC/mouzjl1/FjOJ1eHKeV2ijv6uZvhW
elejvYPqIuiSl8kuRcox/0aOtPS50osmoqVDFjndpDDxLuVM0NrFKO3oWhX8
7DEnwd9jMU+UcIJMFXV3wXv2XZPaPo9yeuNH0vG0//g37dyE9Lq0claGVt2j
PW1wgNWPBe6060AjFYWIPk42NsLAeMfZRUX96s2tXdXkhF5p8h066klj1ZPX
OZEUloPhYc887HdIdhbF9qt22K2NG6BA8c69oS/O1zHTrkYQEHdq+dbArFe3
lyYNgHfOwDdMV10g4Cl2SkuwvfXxxN6wWVNaoRkQVa1QwObjIbIjCYtj1Qc0
xJbqOXz+1OBuyXhvoTJfnFgmDtAbceL3jzcPU1qlSdXUQiyKaDKkceLILe3b
cdTynUUD0PTv2NTJmQjvjZ5wej4Y3XK2B4cCoZeiaVE38j2H/HPS8Nd7q6jZ
5Bq6GFZgP2BXb4d1OpmH8+e02xjRBO01C8At84esierjekSGo6RnQwlj1QNY
hkhK/7MD4oDL0NQ2xGWDhJCocxVTYwNeYzei3Y6pEKrfjZxQgE45D5PzIhVH
4MMxzHU2oPPlz9gf5qZ+ziXm3tCEDQ43lfZkAOgWaRKVpdU/oMzErz3PvZyB
c1g639tQ/zcQyZL5KpNghar57IVw+r8eNpv/2cYSNAeEj9KZTQ6YIXHyc0bN
Cp0Wn3/BCSSVK+JveJbAQnKPbvt9tdHgzDTbnl0OYBK0OukB2oLg1kOMvkgt
SXGPOaH39d6zxsbidlFb6uGo/SkyvQl2hVVG++rwalXw8dRuo9BHaVqFuJN5
wn6xUi0f4luFQj9M6PGLQCMtGd1MuYX2iZE0ointnYdDxvzSGkYDbC+Lczll
Dpt+b1Uxgq2qpH7lB741zUyL127o66D34t25XMUZVY05snSXwMa+mzyK5QNf
mIVC2N1NghrKDmG44ahMZZzU/8iVocUwZUT4euwEJRaVDMnt447mENhLlswc
OguWwDTYpFmYRw6SBLtpasAYjgyFOt0N9HBTKMP8AOkcagg+TBTLJilsS83W
FYyLMQhajzbYxG6GGm2XRFXPzHeNloVC43BaEDF0+xyBGdft4HEpCo3Dp2Yw
oXhoA6Zm0uYsF258XS4rpQC/OkISO0SOtDMkWSflS4Z4DnyA+ibST7b5DHOk
wX9gwn5nXMnigdg4B+IxAOkv7QIcp9apxT3UV4n2l1fVVay7XWRAKPdK0bEW
hANZ31L5elhLhXeDAzrcMpp1XBDib7CwwGyGSn0JerZD3rCzxpJPaAXB3Sj1
32vGbEg9uhP7uxEcmQYi8qYWYPtQOUnRamxJZMu8VzhNb5LKiaUJ8ZFCzcXa
59+VkojvgLtfAC9m5+Zd6Q+/k0rAqOoFkZEb2se0wCqCSrJl9mfgkhjcoiJT
fUMFHdG5tw/1nuoFczZAkD6kelZAkKuf4oGWwkI4L5YHI3B3kT4uruX6kocG
dz45+mIOyc7W+Hx8t89t+0310XmypqIOplMDF+CnqHF39U6cA4neEMb7UGBF
08ALsewUKWnDDwxrA/HexEy1kUNjXXdBZ9WVti+7Abmk9W67spH/CmAn7Wp2
lfpXHPNorJN1n6dINpuZ65Mk3EUYVIRvXSrANHqvpAar3tlORlJx3RJVDOhD
A8KyVValvsQCXCOBOUerbaRJDnRf9bFww/5thG7Onlh29X77MPdWuxUR+Ctn
yQmeu/ying6wy0gUFvYSuWFlzAqO5cVKrrKg77YVVi8Xf6GJ8a9SbjaUubkG
jBH7JIgcDlUZYVJViycQLcqxotVtfnfC4XkQFi0jEI4cmM5CIM61JzMWvV+z
QtYOm3WMulnEZbQbImY6gK9UZ9Tei6+cni1FTXzBNOn2WsL7HDMR7JfMOxb/
j+i3nomNPxXmnVYyywg3YBSqvnNLI30171O5GA5E2wtDK7BbeqPzAp0ChzDJ
+GZiJAR3RFlGJffH7a/kgI0XK3BZJJK9/p8/YTjl6AOMj4pQ3qAFXUINUuyr
YEhFl5dpWSe8RBeFNGn7JFwGXdkXQHaTCqIl+EEI/0bk09Vc0sRhmM3/oNx9
x+ogZ5jsMKdHnxAS8z9pL+4KfdYzjWLme4qPsjqPi8R53Npnzc+88EhQAlOl
+RQUQ0d/WuGC6f5PUuKIigU0wAPuPIpOXTb441L1IGye5orWBovAbmCRbqIC
iEViqOIR73WGCtznQmIFqljBFuSq7MR201orZlyBbSN6ecn0FWs+LK5yJnLx
TcXCYty9x76bjE0Fku1m0ZQ5qPplbwL7IfaHQueWUhZHu5A1/PrlkJaUgHvd
V09INyHmVFYyutA52bpW113Me94CFS32QE2uNCcwiyPr11LDB4FAJnfrVumL
1m4E2+6VXFvJlMLPsBiIUPqUPoAnAVe+ARI3LRblp7b7zESvG2vYjC3gjI9p
0g3hiJiU1pU+GM5Qx/Y19aTmHxW08vDt8QkRSy0GSscqhjKPxVcUZRky2+N+
atuKnamB+hoNWPQOkNO8cwJcjNByVs43o7E0nEJ7HAL5/iXCJfSUn9ObF5MU
6sxyvwFORUiV0NrrlHwQcyeCpsTneXyX2BJeqefeGgLfqUy5qs2dWJ/IAy/a
BzgnCNw+igSweZ4U4ukVw5HOt7yanrwPe5xnt3Y9yfKsWIhU+ZweKRl78/jM
gcOmj2SPiIPw1InmUvZn4Qz2G8AxETefnD8ywMemhma9fqNymJJndG4EMjGW
zBtD69LPqzcR3zOylonmBo+hEIUIHKbgLwMqP78iYSbgPw3lDOqHt+n862g1
xwVEeis/4nC+bpesjFXPUei7PJyRY3lBEswmKNUyg/a/B/Ztz4c3oizinlT6
xmoDUDWgNqpDtVWNzLQVriYis4IP0X+TIIkIHJOWsRSmkGlkldwBxntg7+i7
DM7PDn3BbuOd+3kU8P4eaYzkuetdHNYA/mWe8PwE5HQOzJWn0QNCgymiSV64
gt1YTXT+GKPl3j43yoiO8cUzFF0zkIvlrKYxO5yJw0ndU0i8qDALh1K7JkC+
Qs6yfGh4iC+AFNcdVoo4eGo2dLX8xy40Jm54CauaMU42IMN7vWi4FmoOKs8f
b1doS6Jp6QD6wM41/6Y6yJ3bC51nUIz7eU4TZXYNBRyVhSB1QVeJeh/WI7fV
gZsL+yBNzUSef80e+4AhiGZDaLKJMQ2EpSOvPkws+1QJkhZo6/1Kp0mfdrpk
ojekBgW62t22r0Uhq2aAYbSgnI39oLivLcgMd3ojOJBWIJm66LP5pgHU+7Zd
OhbNPwVgdvDKp7y8sOYsS/SJMWHKscyKr3rtqJSJ20eAMfGOYfOUpUPzMObk
GvXch+HFh0chEBwMtHvjMkVPCNxEh+i2sp4hlNhA6NaTZu0LwnLOZvQENCGa
zxRarLOakkRvJlMLI0P6Ke1XbZxlRqe2wd6Xs/crBK55HLU/P4lHoGBnUxak
h+W0vj/n74e0eYYXzkJHEhGyBr/tBds+B5hgK8KDsGTw5USvwrxRtNNcbWBY
YrW9CvvVwYflB8PPqkK2sNZf7tKreakGUMcamKoEGdJUYEBEjHPtR7AqZddV
irgpCMr5vavewGdiwJ8PEAqSSYPDJF4Av0iBgT1D7omC45GcAptkacbj0smt
6UmbU0xEA+YfhdZQ47j0AlN+CVwSXtqDVRcaH/wUJ64iZ/jc731H2HrsUbwr
REcEDRNVTYvvskve48CoR2d0+5ANKsRL7vHMJ2JNtzxM23x3ONuBmzkUtfD7
9Kq1jQxqgYsJ3EbHCngk8hA068xhHkFk0wKKudqs0C97XVICA8ERqIGpksJe
6wDKoRjUZYxnW8I3GfBfJVaIX0MWpxfM2Sme5qatW5XD0ws1BjHOqg+dkzQt
HfPfzi4YI1La10RsbUBw5b+POBIkTC2xOJ7ZiVMC7LaZbOz3dhVpw45B33BE
T0/93fcZ0TEZ+cIObHPyfKpu7JwK6qZjZJkVfp8GUyWB5Yby5+wNvvZcAa7m
Plr1T3Bv0L44zdWy4uHSq8x8zI7786sa5qCu9kXnI2veQxw4HjYRMmKrhJej
+mVoWuKby5KkfszeXRpX5hsqoJmAP3jngEvi7P3NkYAU+BQEISfXkc9yzahX
qymd

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe76Vd5iQqdyi2AFm1JixIwg7ek/Sx27dOkiKu6T1Iph3Nde9OgbvbTr3DwsujN8mrM5sgdBuy9Txu1nV0Au1GQTpCAhflODs5v8e1XcIHrffBp3mnnf9UVgNk+nz1qS6iYlDEtc1kr887/VvvzP//hWqLGI83+W3AedjES639j6YFZxORPLjnYPT+rydrJ51TzeB+E2PP/VIfkjm/2UomTrg9tp0P6QlUN3TtAgtEfks+AZKJ2x8h9AvCCr/w4LBT6I+y+ZE8WQnBWPPv5H8UOWAtm7qwiVzR5migMO2nJs6ZEhjbavzTBMZcQBNIHYuYDHyeTZhKOMJEvIMMm4vF0qkXFYLuP/yBkb67hAhQLjOdV+Zp4b7lXS9j8NShFZl1rJhxg8HIPLiqcIrFFhbVTwWkaJRTYJ29YN6DEqhjiQup/YgFYzakvCuCAHLf2URf2hH19eXgtCt5a4etSMlm5MS8Q3Ox7i0MGBUIGt7dui5uL9No8qIlJTvyyc09Uoxu0gFoRzDjXSexcU3HG1jDEGpdOQvvXDHPLjWzFZN5/qX1HAAET/fG0Kd7Z/mnKmpB8hvNDjWFD4tsGB/P93itbEaeQ10Oo9hX3UyGd5IaYUA5K3G6wGXkYigTPglz5cYnc6tm+/An69qp1e2TSUE5ccLLDBRsOK8ohCp7Bs7qdMZRQPxv9ZbMsPBJ6ye7mZ5+t0CwXPqpgF49s4oAL+Fk9t/FhJ2kogEJwLFascV+7tfejHBUNNAY/rthK34cLh2KlRlurQuLXJLXFr2AAmsJT1k"
`endif
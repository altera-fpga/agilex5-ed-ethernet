//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QOpc7tCZ9T3Wtr5lB7KWNQ+sJrUsTcZJAnmuWkKBNl3mLFn6dmMoLgucyO6w
Zs3+eD6vFLCpW6Cn0ua3Jwh2ifIuhDhWGA0IRMViCQVB0qbLnp18ZCsB6NRp
PFsv1GFQHouLW0quVNI0z+MZ+HiKstqODlZs2E4LPJWNhQBFL1JootT+yMSa
Idjs5a8c6eca5zgNANrPsQTEUnCfYBZkODrjLKbegWa2xK+tTqtuSWLwUTbV
DmEZsnaWsosp6Sq74gHpR59qY6ifbRQ1+r6GHji+HSrwDr9OudTYCAlqlha9
DAp+L9HYFDcQiLtDCOEvAy20IP2lng8k5DwymXTMiA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mEiLqBSml7gWDxTFdeKFhITspg5JyVhFgYyT4QO3Ggq3GhbJ05WmSeD/65Pt
IjGIoRZgzfHTJozkCaKlOZYHyLBqwavIG+XvW/SAwW+J0qof+4jaOX6sRRG+
I/J9qwOZT2//0teDXT/ohVfJA61tsWs1m42pZuehV31yUQcLlho9jIIIl571
oT5US6sQ1L92D58PsCXABl6xeG+U3teCrXNEOkD25rRQEm+AF6qslaSAROZv
w0B19s4CUsHW3yIGQRNNmUvEqUSKLpgL0VXTV2AMr2EMdMcieE3Q1F+pa/7E
438AFUqW9kbbK+fhahNKthDOBeXuNdn0gTq+VeuIKA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iZ+44NxrzgTOgJML4fFYL8m29NW7D1q6YgkSFcdMeQLlJyZjpD0meNSpJnsB
jQM1tXgDxojYPfvN4oiazlcVNKZF/2C6md0Ei3nsIqp+/+9KbFzczL/yLd1C
N7q8+aFy3lxRCd/jlgDEu/QyI0/AjWx90+0m7JDuGwnHT14dY+kEoMm4gLbI
Z4m0DmDFDU1g3GRt2ZzU5Pq2eXOMWb6612sOFWDQ8cBP9VyR3VQ6w++eycRZ
O2h2Ri90jhT9hWSVb0oHG7kTwirYSI0ohaOvbb8KkpkCbhVSILIerNJnIIN/
6uMBWpDmAotlDATpi/D7CxTllFOuGKxKJvpF5B3U2A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RI/ebITtceGhcF89CFETJVTUbaN2qJlHNDqrmeL5XEohJhkjucbR3mY+TKut
1O5XVRVBLS3IHRI4ZsSa+sQBDgSP+WpSj1G58a9a26z5GZBAiEwdrvcXTNSR
YaGMTaIUvc/xLw3ls0sfk+HlZSKiLBf1a3vuUN2snin5SbBQlrW+EMe9moVR
fIMY9Mar3IeasxMQrpElY7/l8EYvkMrD1y5U02s2/M55E6AR0RAViC8+33bc
6X2u79z9XjjtVUPOTj+9K4yZF2Duk2ytoimjCRGRQFvA7cvTzeSFMOl7RUgE
OrmjBfKuh3dgx59+t0RbnFbYPS9d2G+8JbLWpb7eMQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
b2a/lymPdzLaRRGcMWWkY47EZpTzGZkDDExP8nZva5suIV4Pzboy+VkKf379
e79Cmqcao0B6uXrsbhL1n1G5SY5vB0ZKkeXO0Y/facKTJY4J2MAflJx1jB9W
sgR5nDtqQwrF5zawZIqOInkKHw2Wk8BtfbJ1VELSaLr0uEAQ9g0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
I2HoEYEu4ZSy3TegOiv7UGTDslhHKniUtVWRuSE4y996pgLrRtkPGLV6IoaY
Rvq73VhQnHNleAjiZu+l7WcZhZUa+8Y5zAnnUDo+OfAhBUTnUr2DXGnqeImK
pJD5DtGF8Jr72lQjZtCFg1E4mhF2VgP8P/OcKjhcZWZyYBAHcQCsa3V8EXiV
uJt2L3r9jiZQeXfAmB3fO4kjiqBnl7guCZ3yfTK6r2QbhtrUX9MQQZVorQfB
J4tEeOyxmdzlTa2QpjtlW4zuZD9+GJ2ckTWV/t7sZhYb3gmHAYGajXRhju60
Ag8wzTjWk2Jcz32GqlrFfj+FotMwhpLpGxZqC5GXltXc8HIljQSu41bfEO7Z
OhIdZxwLr0+t1SoPLdbotI0MwBxYSl3fYFPzcIfdBtDXLuTHf6LMn4VFtpMz
rdjb8u5Try5fqxw5lLOa7R+tRccunJSmjyPIj97x89lFQOGpmyJcsPFxJWqp
4QeM3nt2J9ODpNbJHE3BxdxJYbO59Sc3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OrV26jiXw8tNa4EUHolNP6t0bmpnLwSoixkfDd21MvFjhjc3HyrrtyEtUKB0
L5ZUcAVjqJ3N3mYNyl5kIoswNec7FyC7GmX6phEaPTjG6s3eAh0F8kjbrSDV
CxCHayHtVfciO7tkXGY9+NOyx6m8yTn0yj2/zEVvbzy/eZWNd8s=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WWWDuAe3jyvUZ+pfgGLpeKiQS0Rjx0PKCTPFtRkN/Nzfvq9LAwjy5mV5C4D7
ecfWsek6SK/PTOUKEct2oIT1jiOLEmY/oflMdjWS2c7iC5VnuT+UuZyFqJhT
jte1Cz3IJKoktYjBRRmLxqczHXLjAbp/m1u8COB5mIbHqToBYNs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
ssEUz9VWyWXzBdcBNYa//FihUvxlnpiHGNnECvfbk1eEIfRYfgnmOia5p/Gl
kc2GZmJQOVaOkLFreGF45U44766kTabBoQgOWxaJNM8y3SmXdsZdIdZTSI5x
s6c6sXG4K1xalxpAUSDzn5+h4/rMYHUXl5yyt00vywHsT6/yLv6XkqsVIbqt
YZOEKOFS6oCNpiqt4ZWvWSA0tPSCr0oBtEgBzoXng5UMGO7MqSDnX5iOcEf3
aT2wzOnkh9j3WowZte1ZQtyEUC+5O6IVWj392Ur4jM13Rt5ZuFslSOR0jQKM
WDGwaXZTLg8ThLRRy717HtwWcw9dOLnty8bZziaLTpnG6J3SI+LPAZssFZCA
iPp8qbJOL3tS5ZigU0N9vRqMiu49tgtFLBdzXzrSUgQOs6XaVVKPYtojNUDb
R4zY8MZ1gI6tIeeXH3yfl4KlKfAvDEuftOyz8GaQ3jIeOTNCOxHvZNIJBey1
25uNbBmQfa8sMT0pEaSoqfYM9VDwuh1NYZjscJiNu6HumlLTjM8154Xct+uG
DoPgz7W7JznqERTKokvKjxTphAKXlJP6zhsBoTsmoCTDUZGihW6HOJGSX3yn
L5Gmc/CkaFQg/EriTFupl1jBjsT+LxNiyGV1Zh4Z8FZkQL5tYl9Azh7ddtSW
4YI482JrE/8/1w6e8QbCkrTQLdIDp7v0+VXwb1ojdWlu+Ln4YrS11QFJqQd5
V0mDtSpHu5gewlrZwOCnvMMuSLfEIq6w5MP/w6MBoHn5bJuKN/sIaAAdRmXh
jSBUVDbGW9zKE86T89poXxSneoo5Cu/5DVtixrrbdDgJCkJh+/K6HEcisOWG
dDR3+3tijclRy642kjX+h9Qgf+w/pJ3sZR4Yw2qU8XbjZIYsikCNAAUpOrLv
k/xAuYuzQRCQtSQI2Lkpu1fDTwTWD+dFfBqMt2awYakCJjbWZLs6y2k1nP/J
3STADeKoGfESmOdfzn1lyrqPll0aCTHLPjlxdL6lu+vgo1tgX24sJSKyOftW
hOA540XUqMFIGdXsWnFU14ZzvK7oi2KYPPnGivcJz1D1GPbULol9tnNuEbYF
Nu50rfQ49SgFKtxboHIdRxqPP64+l2UzDTdbCiXpe/EKGLCHJuqF4Hr7Uoyl
s4fmPrLrRgl1RePM8SXQtLKMfp6uezSTd6aU/6SRJCr/MATetybf3Jm+Z+i2
f6vzLbYwVM/YZ4WkmaRpA3OFFvvbtrxExABmJqfGIPRFMR1438z8ZuuoLgi9
H4DJuGlfNxmfzRpwo9ZYpHSf0ocBEEDNaSn05UoXXj+Y9mR2jqY+kIHH8Ldw
8i16hD3RPA+y7/PMNV/Lb8Lyuuxs9hyG/uPjlYDn+DxUMcELAX0DsHX4eT0E
11umKIaUWDjjxnpWW8Yx9+m+myRryVHNWqevQmESUXxS6j4cxUnHQ2qP9KpI
RRtRrX6LplL9/6W8WaYrdEP7k1yIOgv02kgQn14XEki+HE3paZFAyhjYKwqm
Ix7dsx9G09w+yFcCeszuXlLW09QkGAKiVUzAV5dMZwwNerhea0IkQ6IaH/sQ
7EPMWMzH/fF7ohBBWtbybvS5HVw/0Njuct3gOWbhN0QnJ3oaY4n0GCAPfJbk
26ee0xERec8+O1a9OOOKlOlcEErxas/wk9r47nwTW7/0H4NFwCiVaog3AA4p
XCiTgf4bb+63Ol+/2gYYrD9k2X1iSjqU4lCLeEhtqbKVc9yOB3PzhPahpvSr
55GeOzTS87jDGW8q9M60KEM+w96QofYMphi6628wUmY/5kToM9uDnIHsboTY
Qi6xd46tv2xuIw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NdOh/z3LGtaoyYmSC+C5BVVnr0UAb1ltTHwAhIFCaqEz6kGoYkY6ediorH+Pkty4P5IckEz08IGB28/SMfP9I/PHMhE9lbJVYr6R4FPCLMzhT91Lo735SBGekk4rkgoebNeUyj8aY48r+doq6izRITr0ceVBf5y4K5Q93CbDlDhY9IWU8HWRKms01EECvSlyhl5r6DrDKQpIJvLOC1oCW6Iw5ooE0PgmnqlRjlCA/epy8iGHyz/JMtOaEEbEp97ctSDBQb7RblPYyd2AWiCGh7cL32j4d6MdMBeO55LwwP+MrstyO0kiTgBHE859+oRSpUc8+s+VqlhZ4UijVZErq7gBO+YysHoVi4EfBLIT2AdrPtk8yN47HpOsOLmpqEKbArsMnKB98jzwuIMJgvi0JvDByEp7TMKYuavK+nk5RqSNSOEXlTmbdx3nBLot+/AJOLwFp/3AwbLDG2o5d1Sy3v/TFPh3EB+TqZHP6Dt/NacQRlA1ssHpDwzs4ZcuB8IkJwRexletCwOR3Uy4C6LjCQ9jJ1Ts/J6gZiZuXsWeRvz72iPqns0zznQHSyaWC7/yd2kY/pQK4jrQp1+btfEHHLt9EwQTPPQQ8rK7cQLOxWfwLrebRpTa4nS4Ou86DrUlTjYjHl9hh6vl8lmVKUdXp5odspMu32joSBDjsKFPWwRm1o6QMnA9VoYGtfdRAOE/LdgSj5GGR9x8GsAbdNcvbl+4Jfk5Owo460W2meG8/h88kmEuF2MwkPnJtm753tYUF/s7HSNJpg8raYIZIdB9qunrN7SADbaPK+Jpld6UZTzh8KtdV7Np/ve/kbtTltpqGJXSHAaOD1s6SVH0yuOUjICSQWHsrBJ8pz0hCbEwshcJB4OWzVQ3N247pxZKKqfIVx88iJZoL3D/exLVo56soO/B/cTJUQ5ksAm5JL16gBRxVcOw5c81xWYDI45j7brS5ftpuD6yEmf0RV4qKeVv1RQhI42NCISx/UJ++tz8RcXgT3QWIBtxjEM+e2ULN2gB"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TApa/Theg7BSBa3wEw6qxzgtFnbeGTidOsnq+q/7M2tCOyQ7UjxrKQ4p0sOm
JBFGovAAdnyviXNH/jTQjuWhc3r3OddbJRHNuMw91XDloAROEaIYjf3O/5xH
P1nbk6FPHof58KLgiOzFuOnrrTWB6rbopYNyaFPwzBDjpALOgg2XVkV93RzV
axLXgiTLVK91JYbq16gbZmH551IzQwxk4NGuBmzqMrj3mFM9ve8Vkx+4UrLL
IZ90HYSRtIMnrsMIyzServCes/iHBdKhz8CMbeb5RmtH6rVnt6AL9ySQMD2X
ictI8z+relrVltMLYqe9jsIPCxqfAaYqKxcMjrOAwA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QzUvqGvWW5X4I6JULpTW+AjpSzS1I1cHt+7Jw4nk5wiyh61Lhx/QU5Uepsi3
++Xz99+0vdcPbmOsu98Yzq2kz1kiIY4uTNNAkqJlpxzU4N0euDreOk+rH8As
vUe0L+URrTLn+RUOzLBnJira/BXpdrxZJQNJTDUH2RqBIxVYn6xN7QbYozk/
ksXLpebiVtgdBLq9MIXD8XuhaU2W1JnpwqDlBjI7aE0pCzvISxtYLxA9RgLP
HqUailO1enhiOHGvf2uT4Rg4aPZl/ps6C0UyLem5WSLJtDQFsHzSbjtnxa8k
Xivv+kvyEQ+VSgS+Z/UY8MUJXMM3RTYsNbf9rc4phA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nahISZ5eTS6+Pc26EITH+D2x9ieG0axEPCUgxkXFnx1AMVuYrpO2y0jgDFyp
+fNX/7Q59uy17uoLDedZCxY6KW0w+8DENQkVPuYSlR13Rzjg4ctqOk47nsMe
+vMoE4ij2gCuu1ci0KnyluSDjp+//8GF5y15cONbOtfoZlNxpcRSmOFX6zZV
CRvZsY+aIG8Lcd7Noi0W3Ds2APN4wMLpgB5j+Or8nzXuUHMOhHrOHoon5sUV
L4MpJVDZZ727KW/v581RG4lLdqudBZqy7py0QhzEQK5ECEzWVYbXGzjMUJrG
aMPdc3WCbLtqvmIXmU7E+1x83hrLQTUw/3VLUYyj3Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hsefjK2DcQ5qSATZm9zgFtJ/CRJXf9TpCl5H4Z7ZwTIav1XHGG2OITiQrpMs
0/5cw2hRn3pVvJq3kMp0xZ/4JFNqbOuwaVghJgZOyBa6c891xWq9mR+vy7Yj
gmkoMtCxB7yk2nqvhBnBBKhYukWMjB9MZddQNH/seyDZZtXH4TREDRLy+jPU
VRBsqIIORBS1/UpwU9B/k/xF6PtNpWGkdaFwBOT0XUsKgYQkuAqpxEiQ6cAd
wZ3V+G5wIUYeP/EkxVB985gzk3rVCKq/PkACFvCj8NexdQABO/ESAqWExnix
YCKGn9+EeZUBJbTcRbWe+qLvBpsGfFicTT6uTA+L3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B/dWXha1BlRZp1dkE6Xjz+VTahoUCRwUKR/aqk7IWS3LC46e0p8s5E4zj2d1
RZdPfvQyuLzFxQI14Pomh0TVnVMYudmfh27iFGvXgBp32NeoPsApIcsEH0tA
ILq89o0ulFvCIR4QgJbng539OUJUqISpmtFhAHUg+ZEPObYXe+A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NZg1gZfEPSPYK16E1uv7OsLr4Tna22yD+PMzUGHG1s4VZj8n4b1zVS/84W1w
BcVyNarvsFJhAfc8CCFKIt4cDXViYsNUqp8FvZGzm1QgiO3Q5yvM6ZWlY5ls
iuWGk7mA6zm6tGhIjfg9/taX5WLKxUCYpBdGlU40Q0705sZn46d8ujXuP+YW
on+xFHmW5LH0p2EEhYGSUBJh9ACOvlbNYQTrkaZWce6gcsFQzc2Dw6xCDK0I
Gt8Ox52Mw2Zpcz9+OhMaphCGLtrOGz3VvD4XoT5xm7Byg9IDlBGOV2ASBIwN
SpUI1xLfHq0VmC5wAAlg8hKSDyiyToYT5R2kwuLjE9PMWKIJEJAojn0Oqqsy
ZnPgAKPCp8jeWXGep5iBOznVQpDCIUzP6ngatFJz9xcRhSCbBQgDNASUhTfF
vB+Z1kXDHITKPSR/T+lnOY1+/WBrn69FVLFCmoVAWJqGyaMCTVuW4xdUJQcB
1ZCFsJVzpRvfE2eELvKB1PVZxMe1a8BI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fPvy+xLBxma5wMYjrb2t1dTKX3yO93oa3jboaqYyRLyIiS+6ztENNJMIiXdk
oObyh4rlYYUpqKrG/ykRiRz5tDc0wW7p2IPPnuHFeQV4YAy1D/G3Zn5BMkAh
zRLjiA3Ma1QfgsTUxKPJwTnfAq2HeTt+oKw3On92b95B97c9VBU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dUddJ/k83+WG/7/Q0ngJc8HvP2jieRrqNwv5OzlaOqwHNfZuUTKmF8kfvj+v
91QHUUlXUl101iK2AsJRZ6akjBvjYEUPja8ZQlHXmoEr9T3MzB0W3AXNcRun
wrSMAAx8rE1xaEVAasWvdcAR3fNNNVEGejlGrqYWeiWR8Uxrq10=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3104)
`pragma protect data_block
fdJ1COJYBmGShofwzIuwMU5fcNVU+jtkl8uBw6Vrq36KP5oft8k1IuGCq8Ig
UvtqsOtotfuwvzhk+yRYIUIx66LgPEGvh3+LxcbGgy69gT3AtqTbFstp4wtN
kDPyYRjhx26g8vMtDHn1vgyuEy8g150u2Hfa9Hfx5FcDgM28R1l61XClzLtT
nzIYZsTh9r9eDpDIOTMI8Y442NYR98yZM9XNkdoc9gqvioAfh2Lth9XoMR0P
ttO5Fyk+7tLVgZjphA5r3c9Yn/uGyTrvlkXS8PoAq06y5CGA1DAjxFrTROQk
SWYaZH4MEQUTjDOzAtqTxCpFmM3tLUzLV5L1gptXmG3GCobph/Tf5CtaXN0I
PDilNj5EvfHTZm0Nki5SElbDIK3GZ8w8nVdgjWCzhW2Lk/6VS5uliELfo16T
gMYt7oybR6NBGyhF/gE38w9RgaHMnyirzGTmXrqcztQsTaBYQu0Vyl6wJ494
MTWrYbWVsj5hE5sIVk6E4tDKLmOgR/+f5mx+yH31xAGm97dCkdFdntCxZpUC
D8q8Wsd/WHxsEO1z7NlBmlu+R+LjOE5RfnZ+hNxdzLcrSXn5pjFoWxxhxyqi
TfC6WnoMSP0tcSGWLRRiD5PhwW0UrGZ9G6Ve05YTcpRWRJF5UzUgu7QrZMvZ
Sth4uaC/3k4SvmSE/sdtnyxs/N3VyyYBJlydvVTkg1aqkg3EeHViBDIrllwD
Hoazb4TXHNVpO99e7x3Lx4yrJ2d8tPl8+oUB1XWicxhSoOICJDeedJXFQPvc
QAh7IE4N163mF8Z4zA76AxnKMGr1NWpyDvqM4UGLRX65EJbNPOQy7XkLiQBd
mGHa22buSxTbJThFjc5bchQPhsiZk89vhZ9cdWKDpcPfvUg9RkdgLLU1ggbe
TJBbTSAWFbQ2QQZBsXZYluUoDE8O4oZWiufvcZ51yJdAAACcdALX7vivi/cD
IvH5AS1gTRTkVRNvRPn5va3hkLjSLTJ263VX/12cKuesoQbZjQ91k2b/PO+B
GCJSMNxOCkxOv2zxTpXM1q02Ynj9eXykudR7fjgsEIh/FxI2sujREjPpbEEt
JkS3OUn4SDe+n8gvEn4vHw5/6uii+BLICLDaPfHUYJ2Ag26DpL1HkUUKo3iY
dxENRKPXG3Vdyp5e3wpi8KsubvZ3QrI5DXr/AsvvQZXjYRCflwYo06iulTYX
bOkapi3FBEX7lsfkbdha/hVLXF3S83CFEI/ldU2wk2NFI9pH3JAmllaq1d8K
MoYbPyqztxnUxbIpXsNNnFukqIQWfr75eMADaOiNuLvfh408ayCTN8p/CCTe
llsoOQzu+Z3rSPyWdljyE1SPsjd3iKNH5h4KtXG5m0IEPcW+iZP4LN3uyrRu
GRDYy8VBDRflss9DJfNsPlBsOdXZQ22CkYwmt8IiR03b3cvVuQdxU8yiXYvj
k5lxG5n0e5FP6wcCBZSJKtpwE4aaZ68iUReyxByhuD9KC7Yg/Xo4actuoHE9
CVhsL8wuRu5oSDJHaN9w1Ogs7A+HZdUm2X//jHEZR07wmXa7otCZIdvia+5S
KBYcmGebj5E4J3LU3t5+QvyBJAgOQqw7QlcXJUw/YEs3NAyGXveUyV50egbJ
3cB5r+on6rSWBojgwrRMkstl8zq4CibZj9ceEPKbOHMx1qMRAfWNSSk4R6NH
i8XjXU26+6/NY+t042SLi3DIhx2inHu9fSxDRFxYBk9Lly+g2+q0u0xaI+v4
eG0d/25b3zPFklSsRvaBy26vNPL/ESGyqSt2VLhyQboppnPVtU3Vx3GKqzbL
oQmaBtj57MfaFe24X6eB0xVTObPCWB0k+Lj7FFZyInmMbTJxQ3CJENXXoKg2
xDsxNJVYQECynatGvwXr140kfoNnF2aOXq//c2yDVnbRO7CCLb1ELLO+WlJX
4OlNXR74MwKHNBL6vOfRRm20TU1+wF8aO1gcucGVsLt2BocgsELD6THsufTO
F7qZR6RMZHQvjzpKcfZpnVXl/g9LhLV5LySaslSD4lqMRHVclV/XBKtJDE8z
G2X6VF5li6auw/ZMR0qdLHNRRJNYH2UlUQjR8pZR0Fme6WMBCCJSxMTAshMS
UnVGBCYot+aZwg2GSDQQJxcrTNoccR2dK5wThNVlepj8Xm/iNwnxPg5GXU4i
zzKyNjR2Sk9hXV9bE7t0CGshfDSmlypwl1b1n2Pan8L211fbWmDvVPgQPlKQ
B6AKMDiklmFb14nXtJL7i5qt8lHQvwYL19HTFzRuA4oMCKizGIxkNv6fONk4
03OGkt3dMangdHVl4hjDnGXQlNs5Q71SAzcWMa3pR3RA41C3FMfiFDPgKmoC
ahCCZ3cBY8/iNLgAabQizqw5Q5ufeszxJHOUzSG9bVinUT39W4CYyhvdiEtl
mqSC9jYHDhMZNaVbtpHJusZJtHwgns7AqJ+gajY/EzQB2+ZxB08+4IFXeB3p
LuJ0GlfDSduospMwt9n/HR9T4uHBD1aHY1Ihu//XJ4FYzxuhjuCsl90A8Go7
B6Bs9jK8K8xOiKLRVugctsOjUWWxDoe/4bAUre5QEytzjNGa7lW8jkVs/Ob4
1H+4+sGMRQ8jMP6RyjfyTlU1FHLXpm9XZrE6/wUQxxZivNkG+HzHzZoeoixs
0ymJL50S9KODHJCP5Tm+lYYKKJEzQ65nd/4jtDsxilcuSrSy2iytxIpzBlRY
79RGDFmfuSyU89SzCipDZpOCaExrTU7C5OCF9PV2fac1CgxWZ3arvc1ls8dY
5V3cKDW1n7GKzciefzjfvpTpL9N3kdxFPFzZoB1PaSlFosLkJgGL7BEPiQuW
VCwUAQgJNP3Myrtpril0hqiRTxEly+IOoc9erZHcXPULQRMgA9+j+vMlcWlZ
CTr48qVY+hikfg6JSyNGZbzRZc7ctDa9vMn/RVGgV8lexmUTglQ10Nt1GzqM
cx0iLYBVqdNP/JsKN36FgFPacJet/9QNK2qpaP1SIB+ONqR2jAZIWAt8ybqU
ZfNfKSIRo63xRe/qaCy0JO/qzfSDHmy3HDl+ETxP9AbQn5ZKRjk231iVcxs9
ekoIrQZwRVu32P/1DW8RGRvMdV0NIWGOoNGVNwCg6Mo7LLvDfnKgT3fv1qjN
FHrFDDRDq/voyR6GYKaGyBW95L1QWWcCW1WCA5oenQ54SKa5lQcCjqmmU2Q0
xOBym+Bu3F3LB7SM9VZHRhXsTYfIvNbKQ78zXLc/Ml5oJqz8MNmWU/dsY5iT
56X1u+hJI45+Kdz6aC4epRy1pmKEFd2L64Mmzp/5YbxtUawG6PDmOwebmzA4
iiggfpATfpM/ZSnDMqP/23gA3t4RCqanUthQHmaDOPx6PSlaseMdfyuBpLr5
dH7f32RtKd4Jcu463pIv+hsxzbXT0qh7JnXvHh/nneMkDIjlnPl8VMB0t94h
aqG1/jwfaJ94cddfy1ZR4L4y+1fQH/CB8gV3rlqMDyljV4Lqs/YE2AZ4LsPE
2I7dZqhovetmLwYFtZkMqhfiX8JfbXXwaq9yRi/nzL2wFeuxvL6o74XDusDD
LNoMLaygBDCEe87jrkVgskvAr3IibucEhJvXW1UHaXO4n7u6aFYTGlvY/hJ7
c9e/G+94WIP5VulizGVytNFs1vNewsJERnH3VlFcOAj9BCcQmysgvB/tssQL
ncBTpReQ7T6hk7q28k5Ie4YmL2rvJFrk+faYWe5zNdQ0GZSyPhZU3QUlpepz
WBg6ZRO1j7hrvHU1FFFj2Vi2KZZaUQ3dwv4VZIQOReZcri+EA7j8xQwRJpgP
8cL2BEXIrW6jMIrZ2G00eRbdw8kUT1faLhVb1i0b4hmnpj/O/a/oz6mPWONV
mYg5BcWhYcpVWRXHU8qqXtNeuI2jDXJewC4dgT33397Nr/tBUYGmw4vNweAu
rlLpUam1Hg0YmuC4kU4G7Tgp7cK9jfaDThpcKsfVPZPwbZpzHF4JtXmTlebH
+FQCFVOpSMEGsEZQiPX0uDtrjWkSHkHXMxgGBqvO1dob/O0Fj5ybVfp9MFVQ
/TmTU4lJwpXHs/y03ygGE0s+zBIpTbHWhoYSMWbeOKAPTszTOFCHBuB9YAWW
+E7Q5bSnqgZ7n2lo88ZX/ncCCyeonNRf7UL63+fgrEavt5isVihYKQWL7pk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI1C+7YQ6FpNX3NaMKX5RDy36gcIuFzPR85Ij5JhRxZo6hxd3P3tRvk+qrhUpZdgoecf1rU/GEwQm9mmEf058ieWX+3k8YwqUdbnmDkqEZsWOome6GlRvqfqVeCfoJnohenY59eXmpPjNmHpDGS8vjseaX1QgAeX4IJgQT5Shewr+a9yL2EHzcDBgkf24parSDDpcgUL2oI4Gp/biy3Fn6TT266mvn/r8PG4AvS6Lt13BfFpgi3FcyP4aSZRpIS/XqMH/81k4bn/DQWRPuOTyGH5/6JwCVyuBgVEQMvm+rbvmQfczavbJhpe99Nz3p81csJUoroj16uvm+QqULbTiapstfOJRd/Dm610EIcR3Y9nAFru1J4khx3GhS1OoupviPUp5KcIVplWe/pN4bXXhyn7xYDGqdQteGC24LZ66tAFAUV01Ip4pLhR2a/n6NWtupOy4R0ncB0qV/7ea3fVXss55WfzMel/+qsNOA6RDnq7xog3jKm1YDd4k5ikHdTh3RZlc90CjkJYhxJA79mWLReN37TiDEKQ7Hogr5BBC/qwtsUnHv0n8j3aHoaXuLpk0uKq5aBmEoEKH43gSX0ZkaQABIgKJ0x2Xqc2corkEiU6U6hYF1OivkarB8tMJc5XudThAezhwgCS5WkTgLlVIhEbc8fKThskLOHLvzAV3KLQg7Qtyn6WZSqG/iYxC/6tv/wS0omXME686l2qUTVXz7oeVi60+G+dzqvNSeZJKCK6GwMkc2u+gvKCCzNYbnHMZEw3SMfHxodkZ71Di+sDKj8T"
`endif
//Class : sfp_registry_component
//
class sfp_registry_component extends uvm_component;
   `uvm_component_utils(sfp_registry_component)

   uvm_analysis_imp#(sfp_slave_seq_item, sfp_registry_component) item_collected_export;

   //Associative array for Register component
   logic [7:0] sfp_registry_lo_pg0[int];
   logic [7:0] sfp_registry_up_pg2[int];
   logic [7:0] sfp_registry_up_pg3[int];
   logic [7:0] sfp_registry_up_pg20[int];
   logic [7:0] sfp_registry_up_pg21[int];
   logic [31:0] address;
   bit [31:0] addr_count;
   bit [3:0] en_pg;
   bit [7:0] pg_nxt;
   bit config_rand;
   bit count;
   //Port: SFP data_in_port
   
   //Variables used to send to SB
   logic [31:0] data_to_sb;
   bit set_data_for_sb;
   bit data_read_by_sb;
   int address;
 
   function new(string name, uvm_component parent);
      super.new(name, parent);
      item_collected_export = new("item_collected_export", this);
   endfunction: new

   virtual task run_phase(uvm_phase phase);
     super.run_phase(phase);
       init_array();
   endtask: run_phase
 
   function write(sfp_slave_seq_item pkt);
      sfp_slave_seq_item _pkt;
      $cast(_pkt, pkt.clone());
      _pkt.print();
      if(_pkt.sfp_slv_pkt_type == SFP_SLV_WRITE)begin  //write operation
        update_registry(_pkt);
      end
   endfunction: write

   function init_array();
       `uvm_info("sfp_registry_component", $sformatf("Value of Config rand bit for SFP registry component : Config Rand : %h", config_rand), UVM_LOW);
     for(int i='h00;i< 'h120;i=i+'h1) begin
       sfp_registry_lo_pg0[i] = $urandom;
       sfp_registry_up_pg2[i] = $urandom;
       sfp_registry_up_pg3[i] = $urandom;
       sfp_registry_up_pg20[i] = $urandom;
       sfp_registry_up_pg21[i] = $urandom;
     end
   endfunction: init_array
  
   virtual function update_registry(sfp_slave_seq_item sfp_pkt);
  
    //if ( sfp_pkt.address == 'hfc && sfp_pkt.byteenable == 'hf && sfp_pkt.write =='h1)
    `uvm_info("sfp_registry_component",
              $sformatf("addr is %d, byte enable is %d  and write is %d and wdata is %h",
                        sfp_pkt.address,sfp_pkt.byteenable,sfp_pkt.write,sfp_pkt.writedata),
              UVM_LOW);
    if ( sfp_pkt.address == 'h7c && sfp_pkt.byteenable =='hf &&  sfp_pkt.write =='h1) begin
     case(sfp_pkt.writedata) //check the data bits value
        32'h0000_0000: en_pg = 'h1;
        32'h0200_0000: en_pg = 'h2;
        32'h0300_0000: en_pg = 'h3;
        32'h2000_0000: en_pg = 'h4;
        32'h2100_0000: en_pg = 'h5;
     endcase
    end

    if ( (sfp_pkt.address >= 'h0 && sfp_pkt.address <= 'h7c ) || en_pg == 1'b1) begin //------Lower page00 memory
     if(sfp_pkt.sfp_slv_pkt_type == SFP_SLV_WRITE)begin  //write operation
       case(sfp_pkt.byteenable)
         4'b0001:  sfp_registry_lo_pg0[sfp_pkt.address]=sfp_pkt.writedata[7:0];
         4'b0011:  begin 
                    sfp_registry_lo_pg0[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                    sfp_registry_lo_pg0[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                   end
         4'b0111:  begin 
                    sfp_registry_lo_pg0[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                    sfp_registry_lo_pg0[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                    sfp_registry_lo_pg0[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                   end
         4'b1111:  begin
                    sfp_registry_lo_pg0[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                    sfp_registry_lo_pg0[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                    sfp_registry_lo_pg0[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                    sfp_registry_lo_pg0[(sfp_pkt.address)+3]=sfp_pkt.writedata[31:24];
                   end
       endcase
       `uvm_info("sfp_reg_component",
                 $sformatf("Data written to SFP register array : Address= 'h%h Data0= 'h%h,Data1 ='h%h Dta2 ='h%h Dta3 ='h%h for sfp_slv_pkt_type %s and byten is %h",
                           sfp_pkt.address,sfp_registry_lo_pg0[sfp_pkt.address],sfp_registry_lo_pg0[(sfp_pkt.address)+1],sfp_registry_lo_pg0[(sfp_pkt.address)+2],
                           sfp_registry_lo_pg0[(sfp_pkt.address)+3],sfp_pkt.sfp_slv_pkt_type,sfp_pkt.byteenable),
                 UVM_LOW); 
      end
    end

    if(en_pg == 'h2) begin
     //fill contents of upper page2 here
     if(sfp_pkt.sfp_slv_pkt_type == SFP_SLV_WRITE)begin  //write operation
     case(sfp_pkt.byteenable)
       4'b0001:  sfp_registry_up_pg2[sfp_pkt.address]=sfp_pkt.writedata[7:0];
       4'b0011:  begin 
                  sfp_registry_up_pg2[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg2[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                 end
       4'b0111:  begin 
                  sfp_registry_up_pg2[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg2[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg2[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                 end
       4'b1111:  begin
                  sfp_registry_up_pg2[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg2[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg2[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                  sfp_registry_up_pg2[(sfp_pkt.address)+3]=sfp_pkt.writedata[31:24];
                 end
     endcase
    `uvm_info("sfp_reg_component", $sformatf("Data written to SFP register array : Address= 'h%h Data0= 'h%h,Data1 ='h%h Dta2 ='h%h Dta3 ='h%h for sfp_slv_pkt_type %s and byten is %h",
                     sfp_pkt.address,sfp_registry_up_pg2[sfp_pkt.address],sfp_registry_up_pg2[(sfp_pkt.address)+1],sfp_registry_up_pg2[(sfp_pkt.address)+2],sfp_registry_up_pg2[(sfp_pkt.address)+3],sfp_pkt.sfp_slv_pkt_type,sfp_pkt.byteenable), UVM_LOW); 
    end
    end
    if(en_pg == 'h3) begin
     //fill contents of upper page3 here
     if(sfp_pkt.sfp_slv_pkt_type == SFP_SLV_WRITE)begin  //write operation
     case(sfp_pkt.byteenable)
       4'b0001:  sfp_registry_up_pg3[sfp_pkt.address]=sfp_pkt.writedata[7:0];
       4'b0011:  begin 
                  sfp_registry_up_pg3[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg3[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                 end
       4'b0111:  begin 
                  sfp_registry_up_pg3[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg3[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg3[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                 end
       4'b1111:  begin
                  sfp_registry_up_pg3[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg3[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg3[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                  sfp_registry_up_pg3[(sfp_pkt.address)+3]=sfp_pkt.writedata[31:24];
                 end
     endcase
    `uvm_info("sfp_reg_component", $sformatf("Data written to SFP register array : Address= 'h%h Data0= 'h%h,Data1 ='h%h Dta2 ='h%h Dta3 ='h%h for sfp_slv_pkt_type %s and byten is %h",
                     sfp_pkt.address,sfp_registry_up_pg3[sfp_pkt.address],sfp_registry_up_pg3[(sfp_pkt.address)+1],sfp_registry_up_pg3[(sfp_pkt.address)+2],sfp_registry_up_pg3[(sfp_pkt.address)+3],sfp_pkt.sfp_slv_pkt_type,sfp_pkt.byteenable), UVM_LOW); 
    end
    end
    if(en_pg == 'h4) begin
     //fill contents of upper page20 here
     if(sfp_pkt.sfp_slv_pkt_type == SFP_SLV_WRITE)begin  //write operation
     case(sfp_pkt.byteenable)
       4'b0001:  sfp_registry_up_pg20[sfp_pkt.address]=sfp_pkt.writedata[7:0];
       4'b0011:  begin 
                  sfp_registry_up_pg20[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg20[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                 end
       4'b0111:  begin 
                  sfp_registry_up_pg20[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg20[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg20[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                 end
       4'b1111:  begin
                  sfp_registry_up_pg20[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg20[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg20[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                  sfp_registry_up_pg20[(sfp_pkt.address)+3]=sfp_pkt.writedata[31:24];
                 end
     endcase
    `uvm_info("sfp_reg_component", $sformatf("Data written to SFP register array : Address= 'h%h Data0= 'h%h,Data1 ='h%h Dta2 ='h%h Dta3 ='h%h for sfp_slv_pkt_type %s and byten is %h",
                     sfp_pkt.address,sfp_registry_up_pg20[sfp_pkt.address],sfp_registry_up_pg20[(sfp_pkt.address)+1],sfp_registry_up_pg20[(sfp_pkt.address)+2],sfp_registry_up_pg20[(sfp_pkt.address)+3],sfp_pkt.sfp_slv_pkt_type,sfp_pkt.byteenable), UVM_LOW); 
    end
    end
    if(en_pg == 'h5) begin
     //fill contents of upper page21 here
     if(sfp_pkt.sfp_slv_pkt_type == SFP_SLV_WRITE)begin  //write operation
     case(sfp_pkt.byteenable)
       4'b0001:  sfp_registry_up_pg21[sfp_pkt.address]=sfp_pkt.writedata[7:0];
       4'b0011:  begin 
                  sfp_registry_up_pg21[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg21[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                 end
       4'b0111:  begin 
                  sfp_registry_up_pg21[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg21[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg21[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                 end
       4'b1111:  begin
                  sfp_registry_up_pg21[sfp_pkt.address]=sfp_pkt.writedata[7:0];
                  sfp_registry_up_pg21[(sfp_pkt.address)+1]=sfp_pkt.writedata[15:8];
                  sfp_registry_up_pg21[(sfp_pkt.address)+2]=sfp_pkt.writedata[23:16];
                  sfp_registry_up_pg21[(sfp_pkt.address)+3]=sfp_pkt.writedata[31:24];
                 end
     endcase
    `uvm_info("sfp_reg_component", $sformatf("Data written to SFP register array : Address= 'h%h Data0= 'h%h,Data1 ='h%h Dta2 ='h%h Dta3 ='h%h for sfp_slv_pkt_type %s and byten is %h",
                     sfp_pkt.address,sfp_registry_up_pg21[sfp_pkt.address],sfp_registry_up_pg21[(sfp_pkt.address)+1],sfp_registry_up_pg21[(sfp_pkt.address)+2],sfp_registry_up_pg21[(sfp_pkt.address)+3],sfp_pkt.sfp_slv_pkt_type,sfp_pkt.byteenable), UVM_LOW); 
    end
    end

   
  endfunction : update_registry


  //function logic [31:0] get_read_data(int addr,bit read,bit write,bit [7:0] writedata, bit [3:0] byteenable); //TODO
  function logic [31:0] get_read_data(int addr,bit read); 

   // if(addr == 'hfc && byteenable == 'f && writedata == 'h0000_0000 && write ==1) begin
   //     addr_count =0;
   //     pg_nxt =0;
   // end

    if(read ==1)
    begin
     addr_count = addr_count+1;
    end

   `uvm_info(get_type_name(),$sformatf("addr_count is %d,addr is %h,read is %d",addr_count,addr,read),UVM_LOW);

   if (pg_nxt == 0 && addr_count <= 'd256) begin
   `uvm_info(get_type_name(), 
	     $sformatf("Read value  for address is 'h%h ,Data is 'h%h,'h%h,'h%h,'h%h",
	                addr,sfp_registry_lo_pg0[addr],sfp_registry_lo_pg0[addr+1],sfp_registry_lo_pg0[addr+2],sfp_registry_lo_pg0[addr+3]), 
	     UVM_LOW);
     data_to_sb =  {sfp_registry_lo_pg0[addr+3],sfp_registry_lo_pg0[addr+2],sfp_registry_lo_pg0[addr+1],sfp_registry_lo_pg0[addr]};
     `uvm_info(get_type_name(), 
	       $sformatf("The data to send SB is here: %0h And it's address: %0h",data_to_sb,addr), 
	       UVM_LOW);
     if(addr_count == 'd256) begin
       addr_count = 128;
       pg_nxt ='h2;
     end
     set_data_for_sb = set_data_for_sb+1;
     return ({sfp_registry_lo_pg0[addr+3],sfp_registry_lo_pg0[addr+2],sfp_registry_lo_pg0[addr+1],sfp_registry_lo_pg0[addr]});
   end
   else if (pg_nxt == 8'h2 && addr_count<= 'd256) begin
     `uvm_info("sfp_registry_component", $sformatf("Read value  for address is 'h%h ,Data is 'h%h,'h%h,'h%h,'h%h",addr,sfp_registry_up_pg2[addr],sfp_registry_up_pg2[addr+1],sfp_registry_up_pg2[addr+2],sfp_registry_up_pg2[addr+3]), UVM_LOW);
    data_to_sb =  ({sfp_registry_up_pg2[addr+3],sfp_registry_up_pg2[addr+2],sfp_registry_up_pg2[addr+1],sfp_registry_up_pg2[addr]});
     `uvm_info(get_type_name(), 
	       $sformatf("The data to send SB is here: %0h And it's address: %0h",data_to_sb,addr), 
	       UVM_LOW);
    if(addr_count == 'd256) begin
       addr_count = 'd128;
       pg_nxt='h3;
    end
     set_data_for_sb = set_data_for_sb+1;
     return ({sfp_registry_up_pg2[addr+3],sfp_registry_up_pg2[addr+2],sfp_registry_up_pg2[addr+1],sfp_registry_up_pg2[addr]});
   end
   else if ( pg_nxt == 8'h3 && addr_count <= 'd256) begin
   `uvm_info("sfp_registry_component", $sformatf("Read value  for address is 'h%h ,Data is 'h%h,'h%h,'h%h,'h%h",addr,sfp_registry_up_pg3[addr],sfp_registry_up_pg3[addr+1],sfp_registry_up_pg3[addr+2],sfp_registry_up_pg3[addr+3]), UVM_LOW);
   data_to_sb =  ({sfp_registry_up_pg3[addr+3],sfp_registry_up_pg3[addr+2],sfp_registry_up_pg3[addr+1],sfp_registry_up_pg3[addr]});
     `uvm_info(get_type_name(), 
	       $sformatf("The data to send SB is here: %0h And it's address: %0h",data_to_sb,addr), 
	       UVM_LOW);
     if (addr_count =='d256) begin
         addr_count ='d128;
	 pg_nxt ='h20;
     end
     set_data_for_sb = set_data_for_sb+1;
     return ({sfp_registry_up_pg3[addr+3],sfp_registry_up_pg3[addr+2],sfp_registry_up_pg3[addr+1],sfp_registry_up_pg3[addr]});
   end
   else if ( pg_nxt == 8'h20 && addr_count <='d256) begin
   `uvm_info("sfp_registry_component", $sformatf("Read value  for address is 'h%h ,Data is 'h%h,'h%h,'h%h,'h%h",addr,sfp_registry_up_pg20[addr],sfp_registry_up_pg20[addr+1],sfp_registry_up_pg20[addr+2],sfp_registry_up_pg20[addr+3]), UVM_LOW);
   data_to_sb =  ({sfp_registry_up_pg20[addr+3],sfp_registry_up_pg20[addr+2],sfp_registry_up_pg20[addr+1],sfp_registry_up_pg20[addr]});
     `uvm_info(get_type_name(), 
	       $sformatf("The data to send SB is here: %0h And it's address: %0h",data_to_sb,addr), 
	       UVM_LOW);
     if(addr_count =='d256) begin
       addr_count = 'd128;
       pg_nxt ='h21;
     end
     set_data_for_sb = set_data_for_sb+1;
     return ({sfp_registry_up_pg20[addr+3],sfp_registry_up_pg20[addr+2],sfp_registry_up_pg20[addr+1],sfp_registry_up_pg20[addr]});
   end
   else if ( pg_nxt == 8'h21 && addr_count <= 'd256) begin
   `uvm_info("sfp_registry_component", $sformatf("Read value  for address is 'h%h ,Data is 'h%h,'h%h,'h%h,'h%h",addr,sfp_registry_up_pg21[addr],sfp_registry_up_pg21[addr+1],sfp_registry_up_pg21[addr+2],sfp_registry_up_pg21[addr+3]), UVM_LOW);
   data_to_sb =  ({sfp_registry_up_pg21[addr+3],sfp_registry_up_pg21[addr+2],sfp_registry_up_pg21[addr+1],sfp_registry_up_pg21[addr]});
     `uvm_info(get_type_name(), 
	       $sformatf("The data to send SB is here: %0h And it's address: %0h",data_to_sb,addr), 
	       UVM_LOW);
     if(addr_count =='d256) begin
       addr_count = 'd0;
       pg_nxt ='h0;
     end
     set_data_for_sb = set_data_for_sb+1;
     return ({sfp_registry_up_pg21[addr+3],sfp_registry_up_pg21[addr+2],sfp_registry_up_pg21[addr+1],sfp_registry_up_pg21[addr]});
   end
  endfunction : get_read_data

endclass: sfp_registry_component

//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U601Tn/8WewargYNfCtojtks0UTugGYyR12IGyGDVSAp3LpWX11Rf0Wht2kh
pmJjkjM1dBdxjbQDATo1yNsd9JzaexbFyODDTgt9KqpPJ3VtMb4p71YpRq2m
ya6Db4fqWkB7EjssDTF+BRrFN7ix639rc7UW59gk8X5CYhO/2MoUx1WX3RlY
BYL0JUmTxN5TwQmDDmNl0yLSEslRsG7JKhpk7w4W2e9zY4cCYAXMwL7aUDy/
TlnvQaYN5MmVqZe1gbzYEegP/KnsMwIPZ3qmEgnbhJXgbauAfS7CnYe68/l5
nQCUm2ZU73qDSDPlqJ9/RqxmG+OvI0nRUDL6vaLZBw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GxVi0SNlfaDcf9JIrQPq+xqBK4FRDvDG856GTMnTGlr+FiUkFFiJlakZfXqW
6mFgYYgvLqkeI6b+yAH6wLJFk0R9DqHHRyCFLg9HBMcuaGmBmvRgdheb+ixK
svzyhgPXSczEQs+KtOOWrsgeMuCK0pLTAVOr4QFRYfx9UlG724E+813Sw7J2
vrrlAZd8R3OdyTaRPAbuCKIlbLQ2UBLypCXhKTImHx+6zcRDw/WeLz2n8k2e
RYQ83Z4Q8n2r6aeIb7UQPsIfAYc10Qlj5BS/xORMfMnmLezsjctv286VUs7W
v+GL+MjHH1QuDk9SbKTNlv+RiGI8Aue4IqAiMk1dTg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l0S5ERKnjgLZ5rE5z7KJG4F7avcvRuAI2kG+wn1WB3e/PlXU3xmVbRLTcCpx
7icHzimI2HUc8Gq3xs8b827eHPjuBmLt0fpn+Tr+xKqWM7HzV8ATGobCdVxi
8yic6e4GWT+FsZkj3IC6Xtyx3JvJ7zmcfUSAweeaxW0s2f3KtiLAj+Nv4sdu
eXjs/nl2XCL3KAWp7Dwl2Q2upUZEnYZBBZOENeItmojeKjl+5hxBNobuzYl4
/6nmb2GCAsQq4qpwW7B9Z/ociBCWMyTZUS1dpcwg2S2h+G77DNnKUAyz9SmA
1Q2D3mI0BXorVbB32ia91tYaTkFCiItQ7ovGRv5SCQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i54lV2aXXSF3ZsEBKIUbFvD6tcVdfeMKXimpdlhQ2TQSc6MmP59FWnwS7Tfg
dDsOT56TjDmDeQ2SuKgu5C/CRu3BqlftCsXD60iFJ8k5EPCGluSffBHegHF3
hskS48FSTpKEID2hwIrjhOxgO4Ftd+gJFREkllgMADl+J5IltoJO88UimYgu
fpqEC8bHNclfi9K7Nz6SKo5DGeSHuCicTRv2rtUFgb5/RusYjOZUkYM93wuw
Ac0flioXaK/NQthGRSAGdJ9DrzxbavGJpgWhzFCX7HHiXMEQuSyGlreEaoGp
2Ai4osu/6uvv7/SRjV/f/kfDcAZE/uYWuVTUYOnO+g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TOzilrvYTt+JY3QkTfpFqV3PbOohDyWetYYr8KVo2JRMlduwmmZTMM66LODZ
otvOdUbl/SOgu/akJeKlkZ/QgTET82wn6DQtzTq5v3UMbyKkP/Sh9VhVVAti
WM9/xh+5zsDrRjFU7ySVZKKtKIOoGP4+A9xwBxPuFHWJCh0SVy0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YIw0s97MRjrRoZN/SubgaHXO+P2C7F4ztyDm+Af4o/c1FrfZCiWoyhrb290a
BztEXW3stL5UxliaTXb6geUYUQ+jt3dXaSAnB7IT2DpwpSMH0OdN05rHpkor
KA0moQO6feZsE+uZkmgZfyCtPW6KA6nYeqnOTHWc9pwwcn91LVixGqUoRvQD
Y0HDiLES76MxOEBIaC/wmz9kulgkRVRIlQtjyZj4c+p3znpaXb+rR1QnB+bw
hsbbSgQE1B65DWkdkFh0A/euH7GDl5EcktlEmbc+e2Rj2yWlzKAx2vuGHaiv
DWZKSlvUTY4iWBHv5xx9qRm+GgtBFAFCBgx7X6O9GJwVv5OZP/IJ2qMX9wNe
IznZEf0UKPdN3RbaUxEEs4KdT8W03oD52ZH40JCXhlwrDGcKbUIQS9JSr92m
wq0HwvuYsukt+qlEKs6an21wETAOGNh8NeICMgAlO8JQPDUcG4lLJcn3dBl2
nEfO5O48k/zfzDPsmYnN9Yk2qTvKIxqu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
djlRDh4GnUwD5QrNBmdrm5gaEo+D5ZGyU6zlT8HyURtbLCq5uB6EoRCCcVZa
O8YXBfAbHqPN06YCixcBVXcR4yDPcEGLtl8ed5KQQk+14MPdyrAH2yPGzbUD
93t3B9kEFTJyTHSnyxEV+ZxIuAaoPxebgoyfD7vO7t5zz0w7xRk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QzCqpaokbxwC+M7PKaQFLoBZ5zERkqUMsweyFGlVrXNpg4Np2pPUAJ04LcDo
nMFurVy80FtmMAqGqWdoqRBc3ZNK+0AaKn2UU7dHqLiA4WJL81+wtRupg0Oa
Zdlg4BkVT4k4Wbd5cL0ous5m8n2BJwEo/wNQd2CN05Y/t1pjOlE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2496)
`pragma protect data_block
43NuLM1aPefB2sr3iNv1NYVNMLBOwc3wOMkH3Y1UJ61ncVHj2luLusAMOvkH
4kdloNyoZjJW6khq5NPWvH+ZglTACx00wS/hxWEnQw3nnCaufZeQzSNM+ApG
ZtRJkVTtQnpOG/tdfEOYjOUfYbnjissTqWw/yt9XIAgAxuhXZ3NXJXQsMJIq
VU87Qc4iLf+pxFChIQ60//wCjRsXitT6UzZjavbE11sBOTA4n5Akcj8UO5gy
5AR9Vgkr+mFcHRxF5dbh2pIi4vYEpxhmeoh5ZtHHr/amQ97QdeYWYamLidLg
vI5mVNeQ7jm95YORQJPGSFZ5lK2egbp0PPeXoxxBVjByiGuDYo4WRY9vFCHR
pi+hg3MOiZfnoxV1IMBF8O6j+C3PncwJyuIUqYYng3AgJ0zgK9aYJYddPoeh
rI2p8lZ5lHbuOXevYTKxz+JSqFr7rHUrfVx/0LG/gcZGoD6dALb47+66KvjR
2nHVLwRmL4m6y8GZNzkbP4eQUHlD5X2gcC6h1uKkDc6SxoSr2C4hUNj1vhqo
i9nDALSWivvCaaY3Hd6caD9qtbzEFGvNptCZ+hwmwRVpBp1A7HYLGb9Zq7UR
NYSPnxMSFArUALTBfa//E6+syWHsNlft+lgKeik3IqbOd3LbXykKjVFUUp7H
Q36+J1xV40eC8acRFXpg4dTd38kUnwpmxkM2cmhDUhNN9TwQ9WUebmJ2QdY3
t3lUZGFAH2x03MrGrV9+l1gIUd1s5aoQAde21niDUEMnCRrI0fAL8YOWxLrT
RRHH0y+tueMSTz3WmJtF7CtfT/P0y/jopEak0nKyjnH8pukLASxmggU2h36L
x79Uo3maKhiws+tW5jSzM6MJ31yA6olt5awyIJBiBNGtXhjrW2w8fGgvITBp
s7Sybt5N+Ox/ZoBkUYVONzlqb/+S4l+WE3YGuz3WSTZN72vuLU7MOfDHtfV7
xPo8CbT7abcmZXXIcF51akCju1SZizXz7CvB7Md31C4oFFzSLJbu3jIE9lgW
1TAYI4dL8zhq0whBR21Y53ok5QGzlKvknJKTJJhEn7YZ/HROEfe6bmP/068D
XCVSib2LiOqzVw/XHDUQtRsu2l3wkpzQ+7QHw07amt8Ocjkf4xlj5uVYUAcC
DzleN2fBIEnvSrTZTQMU33x9WEwFebfpAaqrKsWe+jFPWf1Glaakebm2tOwD
+vk15kRARWtlrecZEr32hFc//CovWPXl88cAkstFDCRbsp/wPRiJQYRX7R8l
n5nWNIz+208WJEY69QM9HKKXHIhOe1kYn1KFTt3ONYjxsabl/Z2c/4fuzRO9
zNYMRgE39kUasb5lNz2mZFsVn15oBvtHu6A3mBwVXCVIYlhDaEoKQbRR1zc6
WRwujB39bHV3LHe2/yVAuw42QipmZeGsx39Cb8de6/bBM2PUbxiXGh3+RALm
XDaVhpV4CDXWXwmPdiqIwnQaPJWDn2G+ifZYwrK2QjfHBZTY9HploIc40McR
y8xHGKe8QSKgZ10YZ8ksNXHDMhv23MLOK02v7w0vsF9sa2NtDh0DYnqHkyv1
q2PaJTfAC+NeU3VaJwyj/P3k5CZM5kMWC554s74ShyL8nM3/XtWu1zunWr1+
4W1z7y8hNdyzpqyG16uM1PS4vl7Qj+gpdjNdKQ2cDlHG85+I5BuVDnKINURj
1odZ+qDbzD+ROYXBI9xka3iL5wBdawcEnga7/6F6/cbP1VfkmWTMdLs0ssg4
Cb9wtg61AHY9VbQXsggKUEtAojS81MpIyzTl3zvx/sKNSRks3sa4Z+k8nZ/D
ko3/U4xRv2l2QG3VEipot0VrkrZXJp001BExKtfjcF31WhoEvSnUo86qHFnW
UeYpnFFXndNJRLFbi73h1SvQ/KL5O0/dU6DFHyJcMU8UPrIlUy7SYou+C7q+
tyW6DyW0GNZ1TWPQ0tPmye7FA1NUHLfujaSssefREcnHpkZkV115to5hb+sg
zHvKgRiiWzJ7XrTAfw+qLUzkGI4qEz+YtRDIFALCX2H2woW1iLGc6kHae5th
+u2/jek5JFtTKAYBWDALohYLiQCLxn9TEeNuLKasRHst2F8UeK5ueE3B3T/8
CwBKfdQAK3ruUSggzWOmUHzI9TcmsCwFIaLQ/zDGoLi+gLLBg04K9Rs5DbW8
FrtO47ANYGOCawVZqf+j55QAGxG+sK5Lksu2GD1nMMH2Jn6nkR8KuUZiKdpV
G7PfjqtSBu9jBXVxQ4BOktEhnAIIyUrhPL+YzcvTdfPixNLJSMrLKcRLkyuO
DsvA+gXzK8MvkpRqrL8TuoAHmN89JFh7E+ySFM9aGYZJakb1+xt1QAeyDW6E
8lYbyZFT34fLYuxZ7NZQZ9Kj+OF4WXkIxpW9Yk68MRLcC/DfKzX3ZPSyOLMu
SPKJZSBvwx8CZjHx0nHbiaFG5XXPizzfWOhJNoFvL3IFx3Ii2i4dLiNaijbr
1jMFhxgsinOmrXWU5zs6UVjiVwsQdAVlsKZBN/q9LHZa6nOUa0bLqdDqcYAp
DiYQYfB4oV3asS/GBM5OEJ2HCmzVg2uDygF3ui4AbwLTk+/SCxL4lRQAetFG
zlzMT/WDgVZZJsEEMEiQTkxERrgquehlCuUyOsjvN3Peet7+0hGY5BSwNvM4
g1WfN10YxxYcwiAAfKvUTtPSbaM7bQeUUTchTvH9couNa4oDphcFE/QIZP8k
1DyXhgP9nddp+FDKkBtMfq+59Mj9NA8FxHyybMMo0yrIBxwEg7q7fvF4LzFN
x0R/UiTcmDzr30WEvBHF9usaUjcLPzvEBFg7iIY8FO1xOb9z5HjoVQ+ZMG9y
O+jr6ggV22xFnbc7RJkd7+9+50F9Mjb76mXZgIIj0iXt3+MKDGUCJbEJnGDC
9lwOIyytXdjrR8YVh0UQKNTDIc8dWoMM5EkJii7fWHw2Qi2wgoKTDNv+X2PP
TH4jG9EHiLJ88ItfmRYo8Wk65yrQY5oM0OTujrdLuaPZf3DJ9kDlj8q3lKYr
8+5+EGFV5Yj7QkW/fmOWpW6N/RVWcdaihiMHow0+JNdiHcTsOWxoLNL0Zydv
XX47NollIrPAnNGHHnR2oNslNQ6UX7cQCkowbw79F8wOv3U1jr1ltd+AfjnO
KraGpkqckYbtO9yxvdgHkw7P/j6asQebGP1OlDyzBt03w5/oWy09sqoe8aHO
tgqkGcxYvlO/tLYkzEj2z8ey3xvJIJ46t/+tjpMzqpyX2A7iY6ESWH9d6EaM
ukSFEhoaakoUNIOGaNYOWyQ4Ti/1xCCiapOwm5+lyYxIJpLD7pX6U2aQ65Ey
CQ+WVkHsy5DHPeapW0QXJTZ/w0+9

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI3Ld7o1+Q0dTK9DDnmsyNphBVjeBraDGTMXLViCQF/NvBLZU3d/jq/dP7mm5jGD1Ay6dke7MXBJPWEWHtbPx61kjQF7hhyLKkTYNpGqGXYQ4aooahV0iyjLB9MTtTmiobeg7uJjRqOLxhf2ZRZS4sr3gkBazmJ3B4BGpP/8447KGi+eD71kdLtAfBwfrAbO/5ujn5SvqOYgS20d94pbPeajPSyfHJgakKQQEUZyNkx42vv734zrALFfVDDJhxTzKH8tVa5ZY0g04d5f2AGM8H6t7rgHKi6saBHJHwjcfOp6Ez9pBqBxcZxZuvKfifAOotPjmxoj76zJAbcuZiCfaTtSYhwztDwMqRA0XApA7dXylCG4oh05Rzxl1NYrbIXltJEeT36xH1Y/83fTKju6K5MoPBPub8IOwDXFyfI+BeWSzeYqMQUP8zX8JcE3Xed4w6+Ody3zFaKfM8VHsbSG+dbxJwW1deVOM8jvTd22ZTHZrm3K83flvlPeqzMaZBI6SllfaUZsuzEUd4elbfDYHRNjaq3Sgqm9IU9abz5EnH3yoMlZqcK+dHm3HTH612/SbP6vvC+OFuUOQkiEodthsBaK9rOqs9pB4wT03/3g9MEJrPJZ4/SbYFKpoa2SH3tSrB7iwkBbU4tMxbV68ZdIppWYXUVaY4zUVJdOip5ianoHRDOgAbevXJw7YtAyNU1AeydRFcAV9seof+QhG2qR6jCPugpfMKaBuuK80ZzUMdKuAI/1K2dbZ4XZ/cPKLaOrEFAEl4jv8qa47PWd+DumCYMt"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YMaBI5FGgGf0R2JfKp5B2eljchAAJJAKXQO2/fGWPl+6hXUPykcg67oCJSVM
P3kxpxeIAGSN0APleYm2xbgXBWYO6VA1Obg6s54N1GSyQcCNY17m105dJIQK
6MEmXxgVhj72mYUI6pon0R9lHCc1yhPnRCLWarPYq2WwEg1Qq+GPhe6hBwFb
Ok0L/uMYHRs3+VA4G2NkIiLddlSSidKLYZ3stVoly/IMUkgn7g9u6fbrTrOb
47TCgu3oXKumLryO9PqTweVs86SLkb8ohtz16vN1EBA6FSLcpouZshIfSxFG
q4vrMalSu6D+GwYVmWrCS8IvkG3QFqGViX6X3PY0lw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TEDA6GIfgK1IvWHibjNy1r7bVwWwC4IOVL6RG8mtds+MXpV+SAuRnOM3+5XJ
Aqz6lVYd/kFpoAbYkhT5iToZ8JlXrpU8LZIafkER04dngD8c6dcQ9j5GlY+J
+uwiZgHgLU7IggKOAFh8m9NkxWQHC0Gcv97+4hHSfYH8OXsVHuou25Iak6Xm
HEKyh4eVO5bIAFzRq674/j9jjlzA/ujwdiCmGSSgo6c8+52v4JtqRJT/kX1Y
stLXWV1ejcuJC89q0UYM+b+UVXo7G/irtY587AYoCZL1jGWHvbLfU6JDK4M8
xmFZO+mZiT8un8lD+E4a1l4e2tuhXfh8+MbKSHB37Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TsfKHpXhVkxMlAHnHSzjq5IDTjTqkMw4in+uL/pxH3EvrMoDA3uLbuRBeZqg
+18ptZSRUcTkH9ROhTs523gmcoagTL3c6zoXj+3B82unu/e4BsLX55XYyfbF
afWWPtyHZaUj4l2qHJoWk3bP2TEXbd5IyPLtLkGaFaMdAy0HjUw+8XKXn/sj
hLni6LqMxhagq7HeyhS1cozri2gSN2jv7Nye53CisVOKsv/Ny68YW08x9RZV
IZiTowviKmxpsukKiAOFtNdYXq5k+nZnZh29v2xdFhk7CUpvNkG5y7cxtTNJ
85bq5RQmx5iUGKWDHf84NVHlP/Gg0yY/ijJeYqVIDg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bel60ND4L5bO92gRItKKThM6LU7lfL3lfqGzFyrBk2hF1Qu9lH2prBdptE5a
aOnTzcSn7wCF6dkam0x5LMt+aSqIrp8ZOOEMg1wr9MVRaLP0+gY4nrJeu8cb
dgkZBC7rWKYECBLlQv+1y4O4l1QA6rzFQWs+BgsCnU5unlQ3CHBZ9D6ZRDPQ
lqtcv0YTTJiv0nEmgDWzFGisva79x5P1lbZekCsODdM6+RjUQcZfniZyQJzV
mnsWJi8fgHs8f/u+CX4gewK0rpKEjufjvqrt571juiW4IA8iaPExpmPBhFoF
c8ZRGlIGLqJbX7XpFIUldv7F5O2NIfmVX1x0LwVvXg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
skmdFhQt+nP99yHbbSq6MmBy8+i88cIcO8z3c2CYbUCHnDoj5lztMq8XiVfZ
eRNSCKbWg0YCMfQ2mKL6XrnGqTPI7fzYB+gx3Ldg6fRB2lf+ND+ve5d9FJmF
l4HC6l0zCLB5xXro2iJnS1wUjFD62GGBf8BQsh5QJnGe5uUvf30=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
X8bWQ92DGr0GG+bqjZJopvFrtVBOTgyReWZXMDI4Fajxn+jgkxwzhOTQzbgI
YbMhMtl2gSh+vYqPEoUULztZh7XS6vhVae4n/TLZnc8dhB15ej36MZdjfws/
mGiVkqoBsYX3+JxMwdeZ90sl3NmnVZZ7tkE4ul20uCQDjvhOQxoIUkK73qAu
xOoiiZp1GQzBuIKxLLzr7folORZlHVFt19JN0WooBgecozcXybIUjszMAgxx
DPPmtRLcFf4HF0yd9KbvUwd9wdauRk+3DoHBrwlGQ9KWMDS26jcaJxH9++xa
J1ttMBo/STgZ753ejeuyACH3eh+//dJcWVnv3JwbDA8Peu/OZv7nkFs8n724
rZuxj6wi+GjhQllRjseYzl4+1kvRS3oNC5oDHXVCEQi/scNPPz0u8agi7Fzo
1BnQBD57tJn+/8HrgQFACMuYEcajDi+qqXfHqwmNnRcQsCqxoUvkR3BGifLZ
UgpSAMOuTc+FoPmAp0v4NEgw9L6Sjm08


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rG0sE0hW6bWdgbkLgcAbsd3xjAU6v3ElLBtLSfchfGIPDVtPhXHpW9zd611e
H5E4VXm9VsO7S7H1mg9AuPnurifaCtGD5vbSHFM33eQLCPl3uxey2HFY2Cnc
4/7wNzCXV35pMuSXam9LLXG7S1ick8P5xHClC7ejbX/Zlb5Jixk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IJyaTkCWXLZZSApQIZI9CgHueRocVjRl7DQzN10BqiN49+PhkXPwAwvhoEDN
znTAVJ6M4Hw7vzRPu2XUQbp5B3e66gJiUubA89HWA1BAgSdDsJXvq1LGZYWH
TnZHJqmjOXjLJMb0jOHjqAgQvheESNcRu4EndGA/ALTcftJGY5Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7104)
`pragma protect data_block
ePGNTOtad+521pC0ct4OaTkrdxpn8Xu6FYcSIjSfHTjqjCzwxL+Drwvvyd+T
yHysO0SBtrzqThEuYEqdJe2hBhj7XoefMk5Y2EqmuBfFYn9+6geesIKAdIAo
A37aYvXAKpgDkMkxHsmKlr82YVi5bqy3wBXJRNwClv2DginpuESuk64z1Okn
wyXa/uf5MBPBey8emSwHZ+dfY7Nzl5IBZftYD2Jb1+PiqHVdNrFLm++Hz5BG
CfRj2KFfAQbCBVpDQzv76gGBqog1M4xLEIrNPXodckKnjIejjzZ97eLIxMy+
+97AGgUhw0Rd90+gwQVovFISrz4TXVGZ3dI1stGr1b0AyGhX74e55XznforH
5GTfEHtMVOYbyMQro411fdPohxtfdeKVE+9SkTnZOVUFYeBgErkFf4dI4mpV
XUcioIi3Cp2rfFthkEj/dkH6WYRpJpWfRi3/CHx1dPVM5J7wk9Q4j93KxkTM
CoiHE9Pux6HAb1yI3BlqzypY/BHxbkBpTVnL/M5YyQSMyVvylgwYZX/25X/0
q750Sfhq79n6vM+w1DrC+l392wGw5jTkygJfckFFS35eHxaptJvnOe1Yi3Wl
K0TLAmjHQmGd4RkE71TuL+JPRgnElB6Kle0FUFr8j3otz0h+u4qH/c6TTUju
Y4LprimUsj8MdxSvnH7MpuMe56FG+WvREAGWLoeV8diij8UBUVbIRUNsX/Nc
VC5eAYcZlPQCVQMTPbiVLeeB37iH2srN/3nAMPtAnN8QO4wDxFXSumSuWtcr
7Kc1p+jgVHVjP9yxU53Pp5GQW7LfGz7mhmhFOLnAV8pTHqs5BmtjB6qrIIGz
TrEj1HFBNgXYQybRy2zDXMo8NmT0xWJg07Ga10Ouv8K8VwqrOtyYVL/yO947
bRJmB6YEnJMYYqCQJehZ9qlr7WDtvxfv4PikcxR8gKBDs7S3xATjEu41KNbb
aml7R8LVQQIk+vg78EB8MBvZkQTImQwOqObxTwJwE11jV6cWeIIEj7Ss62dJ
PJego8D28Wvp5K3f0YPYPWlIGSKM/jKxe/j7RMn5yvSHUbwqn+/MHbxjvOoA
KuTIK+6DjEB13Ps0vRKETN3Hh8xfglO7gUrlljFXIS/SInl+2ytSjU3Ii594
6s98HGQuYDcLrR7UZxgmYopIz0GHQfwqJ6daEtHCkWknRaGa4Bi9XY6ZRb6b
1M12pVsDdBKB3k204HctleI3cjy3kyGEhTX4at01JMGnLdViFXbYAdTwsHAH
TnWNJ2YfIr8NNhRJoWmD8TZQ/SZEggE5CVoA0s1nJIZmcJKOnUfwghocs4uv
IJGmV0+fgD4vXNRES+0avDQv+vxLOc+NSmB9gBj0wLqJqjkz5Qi5PPR8ggeG
N6X9ExZFKLMYmn7HPyH1jgnWilzPJfvW3QlVnpctw3e7zRXIZu3l0zCTQ7sH
Vv2trOTMKR8Z5vaSFHzB8M0mfVULWDeNwvs0w+YUwd04v85w1UKOvjn+2NAx
XaeOj42bB8BP4NavthXmSh7bXLDbnTwEAhsJKgE/Aaig3FchmsP1Dw0oxvOb
AH8apCp3wWrGNJJkS8W9LBZ+RFr5qEVStmZKhz0S38tm3x0gMrddrHs0RDfc
qD8Fm+GZD5HqjqxP5ND0nnSPhO1tTQ0rjLNVTBqDhqmlmr/jahr9bQjaqNeB
84KZ7l8AY6gnxkhDIvxuYxmV/vaCna9Gln4vBrtCX/pXbCfHAnheS0ULOJv+
dO4T0aCVJpK4LSYWYJa0TBDqAH69nIJqd7Pw24K9Uw0cTZQp9KmqpebRjV4F
20vs2YtltlHhBCwOboVyY471DODLNLK09PwItso9SCIG8P28+Yg0fl7hFOca
cbHw3xd3h372gS5PU4gRyFVjItFHu1H2lF++JZHSrUSESU/UhFpySIdHdrvz
Mqj/aXdB12JzzeqLSYfMIniHRTStKwjxIWIpMEzKrkzZTx+m9SnV3W6GstBa
ngbQRt0T6KGbeXZJOTYDDkeyrFDfrLwJ4z8eDgmlUCCIwKkUZEivlJXpCwls
YH05segIsq1+w+sKj3Fo6QTgSxMXv9fX/G2JWKFde6sOAcTSeOrrc+t4ny8b
vvEa/0hyBusdqLZRFJRN7yAucEdqa1OSqRxBzegAfcUYBC1dspDYYnzntCBQ
vjGkO84qJ8fIKsQEG+QsvRJQlCi/Ae+Noh14zJ4WG/Xw6eNgmNzDOYGEUMsg
8qILN2ioyR0aCDqIny6uhFK9jTHXkkHq6dRwxtQQyFPrDWRZXWa1ZYMGge8F
liH7MLb/JU5cF9std7P0bddbqkFqlwwDNcWMtZ72lyoPvo5UteuckLOIKR+e
fZLDHo0x6I7Trl7FX8m09LQ0zi7mKgd6zl/PlGh+xpVuFxXQjQyXWT3O0i0t
TWiwLKKP8OZAqOkBvIMHA6ZA4Sk+87nz5gaXcdHXgiCXT0EPNiDXfhDEfVwS
/0VB1XfLcNBc1V+U+gMV2ARmknsRszUU4y/YqtXW+PelAI/K+qYeHFow902e
zksWl8q7B9ZW1o1W426nKUV3JHxD4M2usS/SpwCxf5w+tBWE6f++mRKSXfDt
tfcUCn+WhXwV++0n2OmmzZn4Sv4Ha6gsGV6xUp1hdD+QdsZosbPK0oiClcp8
4sX8ydvejN5C7oQqYuxdUoHQvLe/Xfot+kqXokEOSeKthsfSSPo8z8GkO1hm
9v7u9tuqyYiC0gHFPljvlH0P+CQSO7J1LZjPUYSF7pbb7MR/2Nl9AjQaT1EW
fKiYFg+oB7+JkcHta4ARYWLfcmfffjTL0Oqvpcd9WKTuPjf37x2R7YYE+OoK
2U4qT+mAJWNecIUBiWhN5FHSln4/MJCKNODZKiEQCizcNKFRsH4uplr0G853
g6ZJtNBjZDwjdMhw1MQDfxDgDZ7V5GMonOroBZJ6C6UFNDM3XztBny9EIccX
LBuroPL6fPplT7PkLJvZgVv4ormWTTNz0Z1K6mfwObU8eIRmAp9AiHiAFpAp
Qk4tYvNtUdyD31grV7sDYuSC7e0flYcRb/iLeabfAO+P0W2BRKacJLeXTOXd
NiH/K7uw2xpdeuhnI8NmIY/+6cmkXZSwEgG6JXXgLuA6Vs9NCl+ST5+lDxIp
saW99YX4z4N5VnpWa/yZFjaqXjYBi6tZAdpkZs2w6Md+3j6AvSS9KAkUVKkA
PPc3A1CHNUclq8EaxgCI3X0C3xZiqqGnT8/y2sjfDGymWytzkl3HwU59NlMs
tM3AiTaj/aWl+1xZAc8SDmGyStGc5q7mO5op10NGl80KAfSq7oqjnGqxvR6x
els31pMSN5fYWoxJuLRYPunAfFdEpFQgKZkdx0HX5QNwhyM1x2Vw1N/xf4IR
POWqqbTiEtbr2wP3p4ujQa2I0bkSUt318Ab+wnJE7oEISqvBdQAiOw6e2VkV
wwNeQ5IlTUDf0TWr5FrzfEC8abcm60xZ5p6etVsFhmwi7H2ah5Nj4IRDVnvw
V5tNu9NDvAIJnb9IFuIE//qchObGTOe6cAsrKhJP24kMoK4++3/i3FfzVSVb
x7Nj5UyDXLFomsg6Rjv95VOMHUB3Kqrg+B0e2IOHEEB8O1P+Of5ZvROeGEb8
BfAPFkgFJ1ZwjxZBc3Dfaa/MBC6z5OnoEkKhQowoyX4lQN248B8eII1ztE/w
NHPVC+/1rOYUW69LmVmquHDGkzEY+BnRlI0aSaIRhXjWSbvXJtIcLpJ2sHil
hNdYghSMyDBt52a8k1pz0iKBSofe5yEh0DStmS6RLL0nYj750XtK07fH87p1
s4Bk6ppp8SNaHt13D63NF6zfLeMEuC+XeYBMW++Jj/rc6+dz7zaUXgmTRjQf
0mxenLxkngcmYrj7iDA5VKBheQmUTR1oIXCNWHsEeaH6A5zIozHTe9kBTD7+
1wHidn/OWTuG2IDGpuw7nF3hIUtlKhDlLJceRljni5hoN8lOuZylBzy+R7Go
y+KNC/yIqQkEppvA0Wy7XlI8h3NS5aFrONguc5jd9KZ4Mv0VIrbhv5JOnbm2
DpMVdjMoPEXCTXBkvv/f3QsrtUUhtyhJXNFQFxusg56fHVcET3eLgbqklHxo
Zqjyk9TvkdDVKGbJzAlVbrWYOO42h4gPltqkYTvBHMSTaSwGQiATTNBsd3H4
KvCx3sxfmL3vq9q6vxfYH+iteGXM/4S2+9j8UdRxuy8jaFSWAxkLYbRt3Txe
UKkq4QWLPh2LZjupGJXZW9sd2NzPc3gs6eToAVcWaQep8PzzS/FEL3G3LVcz
hDxnTKP3yF2NViqyBXbOERd70w9zxi1tCmgWXtypv4Lp/G3XdUKQ5msN/Rpf
cMPS2vvXjoISK96//eV7EiABQrtzBsQgwmCrYzKllwzYBEsBsqcRIJeOn9HY
/ReSV+lSReF79uLjA83o9GJmiH3hV4khKyhmg7bPOTa4ZAmX+B4c9zWf3/0p
QWn3uKCWA8jV7qGDl5iHVXjLRAFn6gQGy+gO3yTaeA+fuognAKYpxLyeXZX0
7gsdbm/IW+bgcQbpm+XXRzWOfPLDBLJIwLVYW/jLEez7xPVbyXZ/uhi9FPMx
oiMYF8J1FQNEWPNImyQIaasRHlIeh5JYLmDmEZ5VQ6l6DF2z/shfL6hrr1oB
j1WhmHwwgSjKEcfxRYVedVekWSZAbNv0E7MgSKCRww9LRaC9vmCvoEqYNCmw
FqF3/9HaO3hZBlUyAq5MO+d7EpaFadcdWUb8GJgcpE8UtzvkGxBDFnCwZT+B
Yfd+vBLlmcFQ1k6g1BMN/5c/BS/Xc5oMPw32rrImesQZthYX+Ox+G/q6Lt1Z
DiF7qHzbtB9BGUP8sBBKi/4BKAA2Svc3aIBDIEqAvOMX+d3oS6GxTasd3Gck
l8/T6kdh9j6/6dkD0xsiJCtkL8BN3rz90n/+KNSSYGnO9osgyb07BTpNzkvX
q8g/o9cnQCoE/4y8yoGgj9gvAV0Bvu5G7BH/77IqHzSN9eXSX7/pFw0kYNR5
MYQAefx20aYI2MwqEOiO60k2a7D7ADvL7JxN9HVRZHQAV2Zl8TnRE5K0m+Pb
7ff+yAMwwNu0jN+rCfV8u8dgGAWeTkTVjj67SDfy3UG+PHv+a0Rd99URorDh
i3E0QhrpbhUrJVX6+jKmEgIW/pNwZE2iWIwsW38jY1MTc71bno4OI4DarmSs
dmmnz/cmgPCDERFYaaZuH84TEU3DEsA/E0Hvxtli59FSrWtcjaixkgKKRNX2
l0N2omg616OKg00O7GFEioUssa3iaHQVaFzsPX+tLtdd1PrdP+0cXFB8PuDp
Ri2DUQqpni127l2kpP60SAG7dijYLiRTp8QXJjh2XuApUbRcPnY1gbZZ0yY0
Ui9cE9iUNkeSXeu6CBiX/0mEHp1ErgZqZRlkqkmiwnX9uWZf5J9JynIm+PV5
B3kiWnuxEpqD73nrDAN2ARIsY3jzbg9G8YedvMLLGe9v7TKzC/2+zmuAW/b9
D5jX2D3rqM05cRvbKcI4l0cxumWzG5iIbjXYEdXqqOPxBPbbSgfc+ffEv/Qk
aZAAvayxWqJ4isbfKHu5q8qT43O38S4u9p2LIaVkhDdkAxjdqhsBdlLJqKz+
A0JJsRfHmxcL4cTmHK1HU3M2BH6zkzgoMEihmYyOoTEchJwC3haePUK9cszU
AyVMYw7He0Txqdc2MpKP1Gt2+QTU1NNJ+Bg7k9rvWGUaWntRVj83iiF7917x
HXwFKhNb4yRf1R7g8C1u9+dJvZWJfmPJ97GUbz0ap5qfj0QvPaKCDtuWYYgO
sVEunTLxMQt5HSS6G7+BSxkF2UXWK8WITn1XoVYgVVWjq2YE3xT3EloDdXzz
IKts3Lwu54EV2kbMSy9fmxLf+wsS2bwI0vR9tFZmg834zIbejJ1yz8BclHW4
Ch+ht6y137KB51I6FL0RhhEerYye6EkaGCFe1Vrp1gvtjiflgzpZsniKLGqS
ofu4RGtQ0uNPbKLq2Y+LlN+boBmiP6HCCnCdl6ZBNrYkov9Cow7andxZvd0D
gd0SJ5YMzgVgU6pOOmk8s1chaMx4GounXrp/FjWla0y6T2/Jyd5g1cYpVYGU
PfJ1WhjrqFAoHO95AkeKts4lalMgzoMbN8h0Ui8zUSXtY4KXI5v1nT8nWq/x
UrCQosfOzV0SzBTECuONarRXEJ4QZLQwWvKn/0SNTDmZJAOBMcKVqr4vp4pL
pb7M+Vq5pyjjRP1JbELwTuFCLF4iHYfxFuuKLSOXuPq6cPrgwlx91QX9SP50
Kg29FIKYnLrLmjuos1i4CIT8apLXYTmrI9xm0kQPL0XipiaYqiVcEnP4OTud
+uMFjXhsRcs6X0ZR28oMQhOkGAfCylhoUMBxWv1lQQfAEyj5O3t+FP9dDcWQ
3TWtP5njEXBiLyfy5YtVV1mRj3DlOsFScX3GvMeE4C2V9m3VCk0vO/6ovxnf
Ke4tAf3nQQZS8vpVYJMyAb0AnzlN/Rn2iIE2mlM8dIqJjvY2ModoZkjdZJDA
T63jWfYlMj6qPMmVQJWGIkYtWBvhcfqL1em0/ryIrFAmaw9RrqplEmkUKaPg
0JNk6qSrqNvzV35SWqjwAGxusbSBmVqdw0adUsYB0jihFnLqn/DLS5LZNg54
kuaSl1vH7WvPcQY6T48L40JTjR/TW3rgIXcoBEU8TGM+XoMg8rDUGmbYPtRz
PMbTdgPwSiNpp185VPFnvT1M1jf4/AUrq2KrTsTn125x3g1mIzRRkW2o4eSP
Bp6i35sJSmDSrvJJVzPoMLrWpIdkX4PPnuJpg9K+KUu6EOMnE8nhP9Hdnch2
M76l4/Zte3Wm5S/aXcMlcyju6QA7TPz4q++9DbjgKkzLWvAPeuRwCT0NAwLW
XHVguwiF40YW69LsAjvAd3TZNZU6JWdG5F+R5CK4vcrjRmpoMKoG352+xayI
uPJmVDRkMao0VrgMjPa4fz0q3OjmRasQZEx+DQ/9wb3ObtoMKr0idPS+mcPZ
vIqfVtIrhy+P/PUgiSMrZRqHmOgPTjxFRiyVBFpt+reVFyaovkc3I3ySmjfK
q7P5IyFmz0Bj4r04w9Q+UmykgaQg7ZNVvJ2b9s7HwNDZxVCkBBfZJLm5QVc3
68ObnGWl0zNwdTRCJq0Ry2VSJYiOiY36vCz7hsy+EjIrs47ylqsYeAOiLNaG
8iX5Jh2ouu2Ex5Ht4CzP4tiJ83iu3CZmNCBYRL0h/PL8RLLtDvRbz2ZSKKyJ
cd/CD06SWV3wc8FTzxllJMJ1KLDp4HenffsIgaEHby6P2SmsHsXVeK1vcLOg
R59xN6gsA0qK4D8cll0c7qiwynJ2boIv9r7/Q1RT4aM31PsVlfIuU9T/rJeA
jQeJouVylLeuWAqBfjFtRIiAEFvrcYcz2mA6uLzp6FA6uWmS2uRZEaZRuiJZ
PaAecH806d8ijUjOOwGU3KukG3qfVhXCH226btwxfNFGVCVtuDciKx/EExdE
9ZhVH6xeE0LGIr8MdYc+GqW7WJ/vc5LwZf8V6zRaiuY7TT14ebec/+t7CBOF
yOQB9/+FRfyUsQWg0lxBd+1g4aHgRezacvvq17wAeovwL6mtMfdKDhkAlLTk
1fN616lDt/k7ZMWTeDx16/dN2hxbRLMFcuB+EouxRXVHgng+jDpBkgA3qegs
JW22sFpE727AI9mhW5MxDQH6rpYLJd9watiz3mxB3w3kupQFvhYy7zkXTOgB
4U2ZU3P3EYZYHhMjDExl0+w8rw2fyfaFQCJ3bA0l7lbOLjmtwrPhHAYnC51G
kPMJCHA9T8qQIllmMUfZKJbOVfcqnzCmsVsRT5p0197jNeMnimZTJku3C2Yw
UTzyoaaIPgp1bl42Y1TOD5zjQAxmr96AWDBOfG8Tdrkd2jc7+98DYtR45z5E
LqyrNi3azIUUpBbCpSijQkJBi/hZk2uPtBwd+FyIqDel/8ZypTaNeLt/2WkI
yo/u1K36P/zvA4c+eujmQgDu+5xQXCeVQ8QQNlqQ70NcOl4kfkQlfxcu70ga
976C8CmjpqMbC1d9B1tbYvCfV+/uspBKxcpq3k+Kf61VIewdF1PXfq56HHsg
HE6jAsLcwmQi5G5H4//dtGKCtMCWdZKvKnNjg4sM5NT9BUcmZL7SJOvOOXGO
N/6TtDrkK5jayZBhdfzADxcIj0Fhh6Tah1Q+y8wqxN5A3kIR8GtpcqMaQ6nC
Pf/2ljXIuBPTgyofXE5xkPY3WyPk0Dg4OmYDMIUmMmZncrkapClAKo8KzNow
W5eiEBwl7dn6iHmK24eb28O5xtw+SW6xHvcRCzpm/NtfjUemeCoZmlrIjiHZ
8oQDoKKilG2bYsRjMotMtjdpY/HeLkty054sfvs+F+yz1zkzzZUotE/+gCOm
pUVluVXutIu/TqrNvKpCR+UCrcYB6Xk1dqxak72zHomxnDDTimuDVPyo1yiC
ciPk0jnZ1lFOgI6Myrx+HDp1nZQ2d4e/i31L8hS/wFoaJeGFhVzePiYp1M/1
f5JoeG7Hf1PLpe6aT7uwT6wehv3mum6mtdZkE1nWhpaMAzk6W28gtbTkDbHs
sh+wVGKjs+8IRueGxT/9KtzvFDSFVUwBFdDuYHASTFgzxzktgx7vwEBhfm/d
nNXUTg5LkS6ujVGd/PB5Cx+z3qPB0pojb9tUmEKwOBxfLLEdSN717Ko6ydFf
VxP6UyMFihG7rxuYv/tIgoLvIV+qWI59LHfGWMhZHf6JpWgUzyNLErSPwJA3
kDzeuvn8xRFtlR/Dvx7arOlWpFq/Y8/uBcdv4Tv1bZeeX03aaKFf/RKPREdA
QCs1o2xu/XvXoop7ba3cw7WkgovCJ/Gs5DMacLPh4pnUCm/gvpLAQTKOPK3E
3deW/NkROgaLpSd+lO/m56tEJv1UiDqenx2ZlxA8gfaw2HTaAX0j8nEHUwfH
0TLoK80tBvkSOi69k3XrTVrFH5j7ocroR6u53jeVYEzldvWF4XSjqgCZMWpa
QbPCtgXtW/PEBsMZsr2WIsv47wMFR6MgwjW1cqBNjkiPP40t+IorscCvJrZZ
kiKq+QkQRxwL38lbZj7KG6Ns32U6bkEDyfu5eQT2vE/JxPq9kJ10/ZG1DCcA
hLSFr0wscZnECCxefCGMsjvrrpnNzy6/7ICMiNHHqEDlddcvc+2ePFHu/0/B
1RESHlQJIirdFDnldfVDXJn2GenDc68tra3dOXQtFg36ckBIwtz++2i/WSPT
W4NspcGZFVzlwjXJzDvplXlPlsUz3gIJpnry5ZbWH4QKYwV2P1ahmWd+GG7P
AzeWATzsUo3C65OWhP6JOr+uT9m20573LtWwHr6kIMQjhbwSvzi/5yEPK38o
BA59nbtdiFIAzQoz18kpWvHsCC+D3rJrSHNn00tJPOJxO6YgyJqzTc7UaTnQ
0/wODoE9GxL6GW34qIjBFuzyaoekUWabqYBlgf3tJAzmbNf6xbxR4LF6oo8/
GkRVtHPT4moZ7F2qxObQdN85StYk9YJqTKxt8WJ5HV4ZSaAo3p5z

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NdOh/z3LGtaoyYmSC+C5BVVnr0UAb1ltTHwAhIFCaqEz6kGoYkY6ediorH+Pkty4P5IckEz08IGB28/SMfP9I/PHMhE9lbJVYr6R4FPCLMzhT91Lo735SBGekk4rkgoebNeUyj8aY48r+doq6izRITr0ceVBf5y4K5Q93CbDlDhY9IWU8HWRKms01EECvSlyhl5r6DrDKQpIJvLOC1oCW6Iw5ooE0PgmnqlRjlCA/erR7CpiTKie0aJlvAPi8PjhmxG/+maFQ4JA9Pgki1pR4AcrRrYPkorndKuR5urPd/7vM33KDBlTMViMyf7X+/q2t0CmYFlDYJoYKxosPizBkoXLxQ69RkQGIYL8GbSnsxhSu6/FRuWSSvRy9CRPSjn+PSflk7A1qPwG1G+HXK4wcrPhL2Bs3fAf9YL5Eur++EeKJkrtNJqRLvfHmFfGnw3wM5gfngtT+dBHYaOcCtKsvePjB/iuzZKWy8uTJCnNxx57TJXEwjBbv7iE6jbFFZRiIw/ZqqezyuZiKK5ntblE2iv2MZ+NZK9Ve8uzk5Ca0Pa3scSx/u5xooTy6V9n7nhp7e3Paaf5muROA459VhmALNlEjFQeeGKK1n5pUPtm0gOaKulskcOlOetptAz9ow9KvYMexgrUKGCg5HApjlZSvjMXgUGnmhyU3CeRXhqrwqp+mwuIYzcmn0itvnIIPlUMJ27Qg7l5MqBlJjDqdycEJq/LCDwpN00J++BgJ/P2037Gq4hInhRNU+QJlaXdnTIantx7a5LeC5W/DT6Xs2oFA2QTyhKQGVBXIE/gD5dFPUunyt6eNZRs3BC0baOfSEHgo1jrCXsEwoKRYcegaPo6FYdLbvS5DuAW1mGcHQ9qJYq4LMDRs1bhVoa8MruwYW1EtLQw2yKfHyhdjHUK7yh9IHyy0M/akLMJE2KVJ4eynxfAzhHkYh+rjuteQahJg2EgaufkZIOeP3zdoJtPCIGKsMuX4IoWi1uoFPqB54lFv4q56jRJ2gRiQPoMVCvmCFpY"
`endif
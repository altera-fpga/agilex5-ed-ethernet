//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zfKRxYgpgJaehAWWCKALHWD/iU9CukqVr76jwe5ZQ0vMhzTGi9gzR+/HtO4M
EY4tGHA984+vGHm+ROk0QEwEKP/bIG4tEZSZSVW4MPbXBt/9YRHsnajU/QXZ
m8PCnlk0I8DdIz8RWyimEWQibdZaZsr/HBXKMWboevjDEhp1m05YWLaAZjU6
hOCqEEkBJI5nsZpfFtZYHFtb3UEwzlKinWKzzLqXkN0tawhpHZCX1qkGatYO
LkrEPntUZkJbKw7LG9D9LRmfukcIRB+A3N+mZs8iayGu1R36OwIIJ41Rn2Mv
Dvv5yQgX+IhNOukRyi89IBNY1OSdMGhkTaVvDUGsLw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c0yR8hB5Lym4yKCW3ZScpmvyPM3MhV+OzNvl34NrhQsWJFla4DBtRDxDgaYQ
ofrhaxrNJEqzb0gkaSGKz8S7/9BcMT0xRKLnCX1qe1xarrEaJKOlGTnhikTl
AeBoMcZseMaUXMQMkQ7dYuIzbSnDwK2Wgz3vCIU3Q/gcUlLCW53nF2e4mqPO
MUG/Ro/u9dqE4xLy3XQnxgJrWxkxXzn2kjgYZmr63N4dFPyj+CIEO3dJldKE
LWJvgjg3kdFqc5IrzNMrDnv0pBZvGwXLvWBujkKvrLDmCkdFsOw0ouDVgVel
WJFITCufPTwUTMX+/QW9vE8P9W0LLaleFDFNunJYEg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F6ujw4ia3Q5AxQIR8JHsquUTQLZDcFjYdFYx/beClx+EBNBnZEI+UraXfeAa
hHRAAG/V2JdAjAH7/zbOTJIDhER520xoPbg6qMRonjw133piS5Br63HT8p0E
hFrPkjA84juAP0rOCvaaYaA7TMqcq+q9mNd2fYLh7LKQV1WoW6bT4W0ZGFy8
ZTs8cEWefilkkKnHESpH5rxPTet8a2dCx5vc0bauhtnnPep0PA5WeplUioGF
rtArMobLbGJTNLTQDKx7EfpMqwFvuCZenLy0K5LAIcnOteG8RolyMfOP663G
IgpKWZ0CZ71q69rvSLsrE1vVDZICkeI7Lk76YhCKLg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ze7IqmkjdM2W4erO1BESG8nPCY8WOMopp9ks82KldZmG7JkAl33VFT0/Q7aL
hcwvaKDjPjeMord7LJuVGO+qjDrTGZJpQ1PPLXzDTT93LvrFhxCuY1ZXZVVw
Y2PoYUSla4e9gR+HUBqOGkBWf6GDg+2zFU3ji+shjwsrfR6LVzgjaNCplHfe
Lg4ZMv3imXaFU/7l/JaaJ1z/8atUDRLAx88VFCjOX5LsX232Rbq/p97WcXzK
GTGL0JFuFsyYhJUoIIxZXkQP5Z/xNgsBhukUG/2Mw9Mq+Q1BQV4uvt4mJ94K
8ST/KUIkbjUyvpMNspLQfmSx5j/2/o98c8hxrAkHdw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
M6ZpjEAj8nDxA+JhtLGHLdtyRPD1HA7S383gWAXjgjv6bgSoruQYLntNm+gH
uFw5sIyOvIJYkq2EcCVYPRVh1qdAaieu/QTa6PAMMvG6CktmOj+bp7Ji8jiJ
j/oNlu186OUC5Rw7E7mWsQ6qSqqUmrsEB/Bu82SFzPDjGb3981s=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pseVo2zXoXrlOkd6hVTLxwz/rcu5kLc1D8h5GI700mDriczfdLDdoZdHhXIZ
CT4lTWIUPFrhurhYM5MJctI/a6GwOBzlyntkgE2l/7vufkVCjeZUHrROiK1m
WVZheelN/JsVS4M2nc6vjGZG/l0fL3kDsMvLbZo6/yUMF18CUZJvpwPIXXQW
GN4VT62DsOOdG/42rs1aWozexdtxecGMkMHXamPhYH3TkDwon8PUXibdhcnL
fKo6i3GH3byuu5VMgFe00YfVeahZW/xUzhVBe7XbUdcvV9ecuiSfT0lIhyHg
lg9YIFi/K+UvPfV0QzTzhQZykN7S92xqolpPvNzOHAu7CQ/C9oTY9TrgXazW
i5MVXZgVFakiYIvCF6nTenvLqM00cdC4BFqNfqb46g42qzzCnp7eosSt9kuk
M/HQxrXoYuH5DYA7Kulv/DChga1cIWPD6ySqao1SyqQUssZ3UzP2YI5MnGJJ
Euv45jITTZjPgcA7TICv1fuChG3Is+nV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mlgswlsAJVbqD8Dzr2BJQFegIadFjJjqbhtivJ+usNTJ0CnR9oFcBW+0y9WP
MqvlobHAlg4h2i9+udataa3GUoqctfW5B8JnsrRHQeOhkOyKANEGP6Rs2vxY
DkNO06nF8/KbrKUyvfhKwGJsQ5C7dG+eca/fBnM72hR0Lxue5Lc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GAKCM57M6dt+1XXR/yrgQlcvn5tY7ud5a5sOl3tEOBabTYGdvyVgNgkbNo6R
EGHmhHsSDiuJgU6hvnhdE0t+632cEDAvmSkEYEnfQetajRAtLkLroJk8lfzj
MaYfeAED1aK57DBei60EYBm6psNGxNSHYJzSGCZfdJiYoLYCP9M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23200)
`pragma protect data_block
jYB/NFymQ8cSE0mSw64065YfDCnkt3YW9zE+Ag2ScLcpB7Mq4Mnr7gr/yOcU
nZjpeSuzlnahjq8vyNNbk51zwuFmQtcjT0xQopsL6EWRkBECce6mcFIgv8Ig
SNyluxN5j93qktfS76qmVb85p8yOXona4sD6rIhMNHrc2sSXEL345LucSW/+
+PiSIYyY25TStuojGWU6AOMjgsJyyFLCWX5mKmojT0mKgOFTvbI6h2+PIT5Y
zK31lTFvNgbiC37R1zHpHPxjE6uI+uIDG4fQvVJKxtsRGdW3NrB5tlseyGBc
yb6LNsSVZVH2+wZEIpNYjXXBKWaU33nG4nwkJ4OTKod42kqVT7rgGQ/DVt8C
B+oBicyLv5drNV1CQpIyo6x1zwJ9x59GfmQHQXjUKFoJOtp4LM1GP/2EWAXv
lJ+lZJPBZcfW7okNDC+KHfLWO58aVYvWihSUXRF/tp112F2CRPrIlBGz4W40
ZyuKoAzo2MvOCltSfAvR+PpzKBsg51uSLEVnUDNfNCRS2NqxzF+HfAFkfVGK
dW2rPRRzyd7gzWtSaeEXvD9V9F/oCrhQYCYP2e1uJsnrW4IbCtT/K+9rUfOv
IA+vhQLizelXVkbaMoKH4vviCDulUFyPd/PHHu6K0wGeMtjzyVOAKodx77yE
zetwUoYPTBcHretRAPbBB3mqdxkS5jFYJsFUaIJ1R7jQKfq5s5UPrqP+vq92
r324yob+daIRVYdQrTijodBT8ketOBX/3+Ci30xuCnyB1Al/4R6bwgiw2KYJ
m+NrIO5Kcuv6sXrnke6Kk7reaYlwaImT8A8GsALpyKlizO28EtJr3Gamz4uQ
/3yMhEeKJvVWBaI9zMFvS6/CavIWuD+bfnmREaHUM5ROrlhS6Z8FiZZisr7T
6wJL8PXzQ63urmx3e+p6vxHvfxyMfU0AGt9N3/nr6MwT6XdqjOjE3I8tei2/
UaPv3H0FdxFYRgeT75WxMp/vc8atdVJOGXkFdXMba/oUt54vK08hQ+fOWAv4
zLyvc/L83WS26ecK6vdunhS+v6nfiCtPJK/W4dVlGxYmDzmI2mvSTh8EWZtd
ks0bOndG7RytO+ylKD5CMjFrcf3x2D7Rf3GcObBDoNHbNAnQkhSDIjbtsu3r
BTpwCoEewMn6adadaknLHvcEP2r7fpbJrcUGuTr4lBkUxFJLsII5ewZ2//YX
ngCoiURUYk+HOF1vV0WhbzfjodnQDPR9FY4VSu9nZqVoPb2g+iwgndhwFJkO
UCdfoKhavSrLUI4g2irrTB8IU+pVaJG0JjkiImPkzhQQePFpGFtNvm1VDjQ9
H3IiqjnnaAQbvyrdWnEEwfXs3M+EKaOqK7ItzmTq/et9d88kwxJKXNqG0B2R
J99b1eZheNgtJtc65NukPxt6/sA/QPw9Hm6Sam3dTUuv9Wm8Y+lKQw0n1A34
cyyEHT3yQ5ZR+KK85PWGqBnNDSnm/5+wlEHIY19LCGYI79DIH3bAlQHmWDfr
I0AVitezsbgaS/tlqtUPfGQOdTFBozDXQxx/kbX/hz0AaQo+RSEhxyoaiygJ
Ev8cUpxbOqPIEqseAXp+xykXQTKQmIPc5e6oZeTKDqao9iqlqhp42ejXREtB
kfi1KOGJKGbXJsfNBieVheHDFHbmfcWX9ztXAteAmYsYm7GhsCDrYgvau/lR
DFfGupdCWAWEvU69EHKi1iQvMkZ2tSpqf56PWTSmkIXkDiu86fpaNgjDUJj2
orVheRzdJ/urfIYJ8b6pnj3Rw864okgZe8BGAHYIfCZbUAfbRGumHwLeb5wj
H3OJOG8J2UKC0KqT55ds/umu6Vwr8cwb3kNASXOvF0PUmC8EYUVHvsuLQCwl
tjt/qB3/GgQsNi6E4PPXafZPsJtzlyVq8Y5q9MaHXQEkH7CrmbWVMZ622Dh5
/vXKFxzTk9KMDGb1WVGWFFsL/Da95xicdCGuJQg5L4eoK0HMwunK7DrBE3VV
BJprkvbOcMZGXYwhdC+Y+IVMLQHZ9vaiRnhbN2T3B/iCU9iIv2ttxml+tSN+
vDOEcAiJySLnBPjn6drFroEo+u/ou2xljWrimFnPRRbnz9BVFU+Gv7SuaEXi
2DlyqflmVHNCqGgexOMAOUbsnywS80B5Uv035ROU8j1XpAQV11Q87jqEEraV
aCL0QuZVDE6Pan/mTx7i88HVbDiYYifQyD7H63+ow+lIAKi4nh3cUGP1qsbC
EDkjv1BnlmCb9QeX/Jc8tJwu+lnSDBaIxDM8OcMKgGBOsconHoJtfy9HtqLt
jWvRsneGSERQZVs1BOSrQNMogag1oQtocZ6l8dy0zzYkFEBCivQ1rboUsOtR
EBi5I+wSLuiyEUpufElQ4fMfdviGHihwKOuitXRExxexKOjnejfSJK7lyVAg
e0NCIJ3CalGskIGXHDpGT+YEW0B8jnkYmLKYGasVxQ0SpTLjjaZoUjoZ2MXj
DFeT0PLqSgZ6VUk7zkmw0jFa4FU7Hz2ffpVqeDN3UvFcseROEHxJGvg1bBr9
hSUZj1Nutoa4zMfGMVJumtxAHqtruGTBdHXUkvs3veUcRUAXUbmxUXFyFV5c
EQVyB3y9++DMN+e1dPDmapv0AyPVly5/vbMkzU7NCHjP7zFwnpP2NFVN8bg8
lKLZLkfcaEgeJuNjBwJzHv0xhQiSYfjIMSSelSVfEUXhDmkc7sapHLKuW15j
AEt7r0W1Inc4/eIHVR23Jk/kSsqWLLjZtOQYB8NDQYRjFzlfBZidXLIQiV8x
FZrIGa8HULeRWZaUOov81X3BbmWqMwwxcqoi/++MmO508gM0OPmn9jVkghh1
fjg6dmMsW3rzCXJUoWdHkUHUTv5GgFWHfYudaFIBp9qpk8GU9YOKEi8ol4hr
T/+N+QBXCXGT69zo2X/CKExrFUTEyXUsLv2Mhx4BNAo1h2ljNR5a8S6KwMZj
y1EDRTGYY2VcQ7fxbu0nAO/XrNT6DTv24y0zefnCXvUydbEZh+UHhrIGPN9d
sco9oAY/0tpSCPtSTNe9he7GdNnXZKoHfjGDpSgHF98nwC/IvhPqMtPYU6FN
/jz2nGrMN5oRcyXGogwHnxeWoE6dUX3e8Ns8NYLBtOJoCJpBgadmyw29d4oh
hD1NBCBzde5qLf3IrHk3EszDYrTcGFExdcp0Nftq2/lkECj8J0H3yPeSJ+Nx
mk6x3QcJCBpJpawq3lkjlv+ONk12HNJ8BNavo2cKHyvJKvBAZ6KvzWhEMpM/
rRJotuz7dMgQNKPLXsgzket+j21VGxj2iVxdBJJpeDmahoDUzNSuXjf+W4JE
nIk/C33fW2YjlG95VNCjEVSaw/vW9a6UYhJeYca2GxWKEjXXBR/b8bjZFsJD
Ny9c9+tIh+dPHvrykR/s9oJ8cTpi1E8cgqM7vbJVYqEGeLn06U+20E1mFGix
C0Mc3eoet3U7ITkWnS+T5MoctUPdfKgyfxs3m2JY42IkhWQKvifSd5Gfk1yp
NGQ+xUbzoyYpC/zbXa/Nd3mewSji+tOhOFCisQaMLvdy121Pi0/7/hp6xHmx
Hn2xQzpg6mchqwVxUlMR6uiHkdlxVzGBbWi6qwx311eEMHo3cBqQSKE9NdeV
yvZk2brGPrWrFEAnpFCGKl8RGz2IGKM9KMnzp8w/nPBUZUV6BU6BCiAwg7oy
4NYMa0bJujrlNmKPKG6eJQL3zP/THAEFyS/jOaqJ2swUrlRRVbjbCk4yHQTz
45Xm7LYAzXupOng2fYMRkjW19exTAGIQsr2ATMs8BZhIsybXslj8JQ2vuJ0t
3yApG06j0OD2VaaUKs0t34fuLNqCK/BajE0k2eTkpxR3S9jzlXAby6OvQIuU
5WXkXM6tXL/k7INDKelH0nhhFtEBDAGTgEBnvtWXHa7asYHe7pZQwN85lSVF
dtRh7HPAWGYQdY2RcmwGkVCmfhA4AWsTCWSRvZkPddnFfO/Ty4AnLkLyIr9T
+8OFk634bflBUpD/tPfEtsNxhDlpS115+vdeqwhx2ccGwhaUrvrXhQPKaXZy
Mr2huDqEsGFWeHkcgSj1N+M8mNSi2IcEZuUZhI1sQQBwEY1IZxalJN6JI8HO
acNXiKggAaqguYEnirpZv4wanjzyGv4/KssT9jnOYWi0a7TuBMq5CBSve+IK
0xIZQyrDJv7CLRTHKhoBrfa48gWDdth/DEt636MIODgmt2hkm8LDkygozQ38
jvycvpXRBSY8G6NXr0Mbpgor3T48v62GzDZPZsR8GqmZn007XlNMjIU+qi1l
1QQU2RlLFSAnfdXfRs/2SrMleXHcEMWUPB0bsMwoIVWNHtdqQbjhglQk56wQ
TicNBpk5xeFi+qCfhF1UBxi/h7QU83D4aujzmO4bSh5Fsn4B9S6zDFU0CJgk
csDTtAI0cDdkuHkgterpS8j0Fl+P8bc7+Alz66epV8FJXUh7UjTkwtrdgrbc
GiIvcK0T824+HbX/FDrx+XjzeWncqgJWyWLfayUNR75cFTYWZkL/p9L6k3rE
ENy76n+ajUJkQQKHJQUleyNsmRQkcSAxXJbczB31wzghfYHaDNnRP3VHCZrE
VrRvqycU9rZ86RPVf3qHNRfDEpTfF+XIKQpvLO/e/Y7dbfkwD7xoF6whMOsB
IDa1j2wxq2igJjwcdrltSutpZaG6t1iBRfLwMK6bACjOLLrL5ElBUboLISHp
o2SRDPOmY2Dh4uexAN4Curco2r50M55pCphF45h2h3h04FBpC33HZab63XTU
aNuiG8pvk6w1aijREMygwt7xGtV/823Dr13q3FU9W0MNFBBSXtmYVMhLhX0t
/dmn2RpZJfmLj4InWgvLn0OaMFueA5plG8qw/qU9ZAne4YCug0lIJJ93JRtX
REsKWp8Aac4eeBaz+TMXY93Qz6kb/fbXmzhhH5EW97cAifRI5s6mrmYHKPxH
6DanLMbIkpgu0nG3d7gFwdWcd9ya1f2csX8Fj/a6pBv/4Aeq8VwAegDA5HTj
WUHFdDW7v1geXxXnmEqjrqU4Cf1C7IR4TE6nck/H1v6r74cPssVfcekUTwRa
6XDjw3DVQqQBkTNt1NJd3VU/DR4RJvXCsPLeaOCNMATMvcUTqD2iK7ZXTUyL
QZ+oBgjlu0vliC5Ka27VJ5ZGxXnqGQ/SrfdWPrpczlLOt0MnzRPdwX1dc54E
ozhqpKez40L3UK1NBH6NwAs+E1AUj6PUdcD+A4wGCwr4CKmJlz42eLY7IgsZ
8HJYi65l+AhIOPDWrhStzA84NYppJMTnQ9gv31ZsVPparLTnYaGCQBAkPHp2
8n/YdeqVhjNBokWHutpMJnuqD7oYZ54ETRwX7vEBs/J4pBTfZaD8ABJRZEFL
yfDTvKzqMrCswXnzZYj6n2QfZOsgIXkFj6ZqcsGRIQUQaZRtu+53puBRILgc
FPOZ3QD5exHuyesCe7NlvqJnDKo2tDp1FGVSE0SFlQRgwQOuCbj9A+naFD/J
BQoRHA7p8ktX8C7mhvZvhnpc/XTKXsRK2yNPM+BCO5i2+pUehpR9X5gqid12
d+RlFYoMyGi1ors6brItOdJZKEQ+9zENs7RhCur/X87dkjY0yXW9nG20Rh0T
ueJ5fy6obQy+Vvbi8F2c661BzCtvrgrTq02DymJzEn2LNNzOywDRgfI8dxo5
GFej4GnxBmF8ykNps7kDp9xcZ46WFEHXuYoXJSfg4wlNTIt6LkKM2veU4YUm
o4av4d2W0oENH/iuYIAlTlYjb/a4wcZEwhTtQoI6BR1nKAg6C/mSMPXwjqdz
Ouk6owSeSYmaHelUi7jm91ZCUFj+HWzaeMm3bIuNkPK9lsnjQ9hCw9xgLv7C
s7b9kwccqlVkVnsmFYnu2/N6lm5Iu0L01h6EMn/qXMw+qYWKhhgjpB0S3D+Y
YRHDdHDSFWHjmHoZlHHZpri7mgaBb6+29r9g36l8wBBBRj1POluDTo1XreKh
6G6iCHcjwHRBLOn++T8iOuE1n21QOihOKsLN9bNzyjQyvFZn+IpJ9hK2y0ip
JiqMZ0pSUqrP7ByuboZ87dVRf9qjjijI11hBEBngIC7lAikk0PMySScsUf1p
RTB42HHZOLUYrVcOaoJJUHNdlu7j8QLz9j3Y49DehIRVGLXMcnKobY/bAgOx
v9t4YdICCQCh/jp+5O35gw/yVpf/Yjc6xLkmJ8odYH90OCj/GkJVRdjJKCKd
ypjdEXqj+aiRx6CYrsrnguslXJnwrqdyStH4VhLMGQkUsSUytVrRWI50RvKB
8QbldZdgdcKMdr3gNqevIt3+wQadpf5apIT2aUFhtyScKp6+eLFmnS8aSPGw
rkWpvF7sOzg9QP9P3OAo+QypFRkx6/3SwqVDDhZsRJMubp1NtE7lWhKa1fFb
FTN0R6vy3HYzQMf0Hi5Xy7/aD6FclG9rpNNXwHp5716AOe3k7xmHmSU+vAIL
+A/1nAm3wcW7Z9UQAX6T58Bu3JWaRlStjAOy4G1Dwjj08upHXQsqegy1bRyg
JoFt10S2yIdSZ30mEhkrCxpY/TtRx87jhNtXO5QeIW19U1UIuPQQFVtlxAG/
cZK+Wh2QR7kuAD1eo1u0wqRIPNl9nDOsw+Cjb6YLSzw2qZOYHnCO306Vynai
a7nZ/TwRpTqsKS5prSMzXNsDc17SSD50DYG5qFpz0bRxlF4Xl0l7kT/XHH/2
StH2NSsmIWgxMY5NZSmkzSTiSFm/nXaBQ52Q8F8NtftNF2kDuEYFcjPipO1x
Jf6T+l3XN1VRGEUbiNwVChIfxZ9vnkrBCcZG/WueAPiqDkqKY7hF7WKwNWcJ
Vv32FmbG3xzTjVyrJdOUdMqMp0tntg8KBA0CWKzPw9Rmogv4H3Zkex74rm2P
eMdtU8TIct3ov4OdIefH5L/b2qaRg1R8Pi27VH7LrJYHhISCROzKxMDnVJuY
JWtH9ZcqklhF5a+uVpfZ39zA2WXn1pnVzRFiI4pViHh883aBchdWXAsAYOnd
pyL7W2eJztLi0N2tki3laOj8jd0ypLKlHwnTnhRdcyBrghdwofkTrU5rawUm
3aRpqDAsHcCj04ha13mjRyUk5DyKehFbQb/8WXI4kl8lgmaa9hW+bE1xk99b
0FNr5fa+Y2/vCT2Gyb5ckWsIMuR/uKnot1rOpJNPUlONkYJh45uHeUzBARfb
adKsCW0o+B6iHEY4ld7mDAGstmBMhkZG4Nu97U2SOKS+n7bH+gEtyVdcXL6P
AmjCCPdpW95IlfMG4MXrMHNfGmsyZfYaAdjhepioeXRkamvLarG9207lEaIm
ENYVonz8tT8kuMoTsQxldEOjqCLCcyHw98/OBkKWmeTZIHiXra0uXhKga7Nu
V3GXCTB5PH871yyXPehn1jT3emuj7lNmCpEpVtWlSDNi8mxeKnRQ2XVUOiZj
03sqNGrmZFUnxiYVXI5/hv5U4Eb9IP6fEfbh5cmdczF/cRpIG9vTWNWHumns
evjHu2TyyxLSm3USjVmec0t5PwYQ0fA7vXTnqv+SQ59BzHy/6QsczugDRVl5
NWI34bdfR6ZY1oUk1JHw6dr/ouHroXaS6LDACIdUPxoh6Ybdpd3NoJtS0aEQ
/KHBrmP+l75p5ZsOiVXLp71Ze6BSFxe1pF26noZVHpGwZ7lb4kf9thyW+VjJ
Cf1RTOCjOEZpzY+YZ16tUsR88hRneTj2p5EsDjiuODW0RzuUQ994yh6LsIDU
Y8ouw+mIUTpSx+bUHHhAA/gwwIooMfCHnfVF/fS2ceySXbPGwANw55DTJ6qH
wG83T6lLf9fUDwoqglbb2DAXHoR8BngJSGXwRewpG9X2ZszsBDGu5h4452p4
4mS1adGYz9TH16/+Jb/kNp9o/ey7xwWDGwvgOxvRRSlhUk8BV0W/S/Ou+2B0
MVeYqD5gyaFmnwRTvKE94DrvyxYg10tZmnIByPqnQ88w4fBWt3+xhTrT7u7X
zZ5iz+XT6alYE2rMPvpY9WXfmqzY9uputJq5G/K7vko73sLv8kbjZZkfZKKH
APjye6FQxrgzna4iHt0YxBXRTShPv8dCwL6Ml9TaLvtoTbGkjxvcXxVkxyZ5
FSuiNokxcrld+9jn5bivxDq+zTcnaSTS+B45xcfZngqc9VbiRJcnbSNT3oQr
zp6bU9XywdCKULq0/lkn+95LTeiIG9kCZ87MAkIciYM2qbW/WyIkI00jCKUT
Ymg9xnELurZ+iRaSFX5GR6zNz0FsABeGW5hZbzrB8ZcT4lMqJWxu9AlfWfqk
WG8L3EcJKbe/i5ZhQ/T0bid35Q2sR8zjNVrp0hmpZXBcadlROXYBD6BxXplw
jY868mnBYXiMNKal+z9W5Rwl3Z2smu9nQ3JrufjmzJbNYgxG8y9hwMR0suW+
Ch1i+AxTV++Nl6zm4Z6iI2xVL+rxKW/TCgq51zayKaFtso2M1cpyVvR8DTFu
XSV0pdH11M+P6YubA6JOTJuwt/syZMYxip7L/ey8ST3QHaISS46IM0fUawt1
K2+5mZ1nd4N5PTkoypS31WF5OOklw37GIMt+xl1hhAcdDRE+dNTmr5HBeUNq
lLe9m6oCu0v7F9jGZ4rcM8cNMTMfpmM7HkO3JL3AAFxT31f26YiavF2BVH3b
xDW6kZZFmuSuE3dy0VxlUOqx5Qvh10bemXdhLTi815ocGkubb9BzP44cciBL
C1fY1llybIiEcveIGJ7zcSF75V1pKXv4AsMrsBoH9oNdneDJ2WwNOuVqOlBR
ydsGsZeucMtAlmU3laqTqjl4TA1ATRjIDSXP2Njy6VzbTEY2zqwPGel7eY5G
ji1qMWBwrzwG7EG+JLgmirosrYcumCh2tU352Kb/oW/cC5TGFXjXGB7c+d+4
3cRustlgt96M+/mddKgGAud7U6IlrngjmMG6kklBgCPB0Y+ghumWxPtSMH+/
LNNLm45KATRx98tSeOyyqa1ygir+iaKGPFcPh0bEHlKU1LokyU3Ym7AHTXZ/
ADcH3G3Gyz2hNygIuziW7IiCPS4YXJhCgCeF0SyD8R5Jv9foMQC6vT4wX4ek
7r8S18A7UNDIm/j2Iul0cDq7967yj3T27BFru8jMWomoSlLtUlxIJ17wBY2p
SfRXkxCdFaSo2yusuRh6TsF3+N4vxx3wmVJicfBQh5UisFz2LjtJhzld2005
lViOCZa9oriWN92UBHxW3dG5wtDgg6LPgZYcx2+lMGQ7PVLzT6z+ixb7+qr+
o7hwr/WaDrgftKH35q1YLIa/Ale/89/hbhJrpTC62NQviQ7DlnKinn0w66F0
lzoKAlIov8y67bUFaZWjynRAVY0LIFWxo2jzMRkm9RHRB31uXk9QgPCMis7w
5gb1APob8uqdzNjColQkn1CJmgKazV4QHer08WgQpUFIwUjl/RatntQZyidO
qZkMVnbDPzCup50DY0RA37LOOCgd8UTLp77xHlD3bInSlLSaqXWzK4tVcfB8
EztIOxt1lkCbzs2duWc9nQsImpjyvqlZGFn3GUO9XRDBtT/kmZiqDejJeOkF
NZV14LVdKCrDqwe6K/Jr/u0jQLm4/N07uaHaFjW0nN/l0Yq4LPN1LS1mDfEq
rl78TRciOg9hHWd5wxrvaSL7SbKJlILu7StePVc2weis/v2DOvVIfWe61oex
+Cj/+KA57VyRkIM/0cRyuI1k9OgTKDMg/A6fB7akl/X7bsb7WGgboAu04+5K
B2sZP4GwDYkSGUXchJ+tbE1FGXOBOS3BOko2BVGwNsHP7qNDioPcKg2Lsxty
zeRSxUS+VIxlV+p4xhPXad/4xfEtOtNPppFWs+qdT+vOHtqHCp42PxVG87eR
i+sf0k8mF+Lk6N7Bt5hW9srs/sM7iiL93TUBVC14eIwx5ETOLm6pHQndZSsM
vy4zWp2/j+irwoozHirtauVCaKy1TV6KQt7Vzzg5Ln6AIouTtwR4f/C3We8f
rMT3cLd0zz5UNVwL6c2X+Cbhe0HOT6yk5K0Mx+qiyx0M8pKZ2+g81GPu+e4D
UvE/17dgJWaHDFQU8PPbnBH4gEJT2FGtH2HQGVd7b91wGRVqYzzKv7iXLQeA
Sfk954OHO+L/qHFZfN13shuX3Qm/S25FW9lt9FuAPdpJlYnhHbF/xg56nrJF
OhTFuOhgEX6Qd7NeCa+2GqkoQRv8W713Qn/AEKMKvwOZxkPLK8etb0GVvPgl
IM5QUfCXyxt90A1xqwSP5l5AB6/GI/wnWk4sAbjfMGk6l4tKbOvyE1x5sC7/
RkT/n9GmAsjduU2qyhobKX7hQGL9WfKPlj7lKytHSKGThSavsqJYF9VsLD93
qAStk6KVMBMr+aRoHq/ifhJdJNI5z5MVLKapi2Vd7ZdTMLMHgghNI6X9Glnc
oi7WiXmVvinRDCSmaun8iPFLdi988BW+NsFccP936TcbMcMUfQu1Jr9v/gmy
/VfJrDnWzt9UKGdP3yEQSyFb5J2Dk+p3yFWvvw2HZU3OuLSb8fMth0pMmpYp
FWl2Zr3j8mx5vROMaLt0al5urGzBs9noB5PK3pyKA4rXMQx1zmUpur7zgEo2
MFEC0Y+Rl33Wu+qgB0mSyflb42ePH0yWnZBWWmSseW5IIZL6G5WhitPXVxxA
8VCA9L2qs2sZUtwLkMUtyHUR5VHyhmIQ7NBikAUdVxTfB+hRWGDxGNpsxmsZ
k9R9sE0YyWN3UduxgPkJ9+xMUT3V16uO9aFI+ob8phu+a9dsUu7YK40tm+zA
YPol3qSCgYr803LT49/JW/ueBpKhCgvqHZYFUXJNNQUe8SZxwrfZeUhG5779
1dnMlpUS+L1vkHBwa9tHRe9RFJz0/oXr59OL9eZX5LC3Dutm6NYqGmNyvb24
xkc/wJWj9F+873s3AreqwsC83SZk3h0HltowOMs754aML2yg6yr3yZS+oRoh
XsIZE8a2l4Y3mKxjMRgg0jPGw3c9eh/RroxfrYFetVV5DX6TUm+P9II6cJln
dTN8AoF/atIZaywhqQ2uLKPfLoIApjm1EqzVUHX1qX4VUmxlcxlwaty1CZJe
NF1kGy9vyMjNqaDFOQW69Ny2VwyZGzrmEVnXu8Kz/lLrdU29TqWbpnZPk7bd
npT7tRKUsVjIkiBcpp8wFk2WUIV5ddol5Rhl/79BcUsHAGjatrHvwEYnsXCQ
SL6o2gD6RJxWLw97gPBawqtQqe/NQv/IdXAeyFLyssttV6BFzG4g99Vwy54q
ID35mYW8iupnV3s9CSiwWLv9kk7QXkNRHzf4AAR8K1oLIkXbUZ7o7QXLkm9v
IsxjcyLZ6Nk57CIjekFxzvja88vIfHs6lhVqGaP9LAM9wWkheKadl0U0sBCg
3lFrrLaXEFuZo9l5SLEOWNElqJ9WNJoZVG6234LE1kl+AuYadwjNQZHKNqRQ
qDf06UVMbXNrws+3uo9fHtZ9O2RC11YUdM8baJ+KEXQD93SruKJrRTzYjNfq
eE8ijQDx+JP6RnowJpQ7/ZJhbo6/QOLV5SXyqplX0pR47UzYPykZZZg0ZfY7
LNc//2ZS/62Gg6/AjZvTLOmTZCTk65kXRdAXt4E+IQK1sQTJbmmeriJHmfbM
OdgmHgug3YrenDZWghXup/7XQzTcUtHa4loq/USvRqzLEa6Q2yWIzuPtBgI9
K2cI+86rcm/B+4XuYP9RLBNcRg7YbDLIERWu4QF5xjqHxCXvIn4XryqT0TGV
IopnBk1o4xnZinby4frQSWc+D8oZuIeCKnuNrwVfjkGioOU2ZlY5XHWTlxZQ
C1+GGPMtQRAmqVRWWZNErPUXmfHi01WYiPgufACijIYlGh5Upa5C1BrrrJlW
8l7hX4Tm3AVATCpmCNMh8qSHt2gOO2/yFySgPwtsLMCBW7Botx3jSa1bLr8W
y0XADBQbRapJTJiXImLhzQobyW3Xrb1dSJ6RPYwnVH+J/dAYMT+Yqzvmpj3/
TGfUwMQbcDT2ShvsyA5bHutr6AgSx8AYVn+ZQSWIPjLyXkCSbmEShvkQzFjx
j5Ws/hZbwQL3fdwzTaNWvCBr6key7tVV0O1jqCYTyxwcmr65zvmt6E+6E04H
4ldWkr4gLlV5jDIUbV1hgI/rDO7dKWSiHRmXaeB5B9LMrrLSLkVYAxkbrsYg
n/efEwxM1AidY/34058fbXYkA0esZ9vj77PDUahFqNCfwyKYdgnDT1F3u2P2
7B9mJx9ZKu21dsirHoM+hoGO1reumivUA8iC6TELE1KB6JNAUgH7rz4oI7Q+
sUucRhME9EIV+XyWKfa+ataicA2ly3MugZwzQII1gDDkqcxc6ctbl9dAXSKp
A0SK9TpZr/0lb/mUV2c6v9a0St6OoKwdRvPHtKhW8je38LxuD0LWl2fA3VwX
Znq7qlLSjIkBXyL3n8n9LmsVbQv4/D18wPuh8P7r/sf4vqVM3U/mTsfQ24xL
+gB4eWnlKEJPMONHnkLZYGmdy0aA5aNJWegvt6oI/GVnDCwIzdtI1RJ6+GPv
58iJ2ZMaopDd1sailP9pUN8+YDes5/kdTnRevhltIYGNCftNDcEjEsicYkPQ
bW3cknkWU9jpJqATLxLn9pmQklpXVGhItnThMSCYHhckC3IIvHphdwVEQKmg
Mu6r9cnTQ5HE19w7mzY4oWwN6Sc7VMKXSpwrn1mxTTTxcJ8sz62hWNomWg7U
FuTA+DLFjE2XonKpwRGj1RtT0gixWsxH0ccxVthaA4MJs2oPXs6XSAz9Y1Qn
1CyzbTP/Ue3Vtql9tjhJf1xKrOL6VjQVWsbFfylmbAhZC60p0AZSUnXeATii
rF3CByiudUMQHZ7bvAGWHoTpAACgd/+UCmFkSVAAI3Fb7L5AY9cQ0/7pNXne
YOwGTyXbIMubsSPerYjDbso4Xj1djrg6lcIjl+TwvhnoNYlX8bbz1A4lL4Lv
WegW7Mzji9YoLi2o9c08slkxy9pIE2MekAuGkrraZYzYEdIpd/R9Qdkjs5Vf
bOzBVBbn1nSwh3uxz2WL/nxz5uVfwjrIE0KwA4f65AwzsxqbMG/kBbG2aCup
P3YtRPLHRmWlCGfxP5mMGDu+1eP8Eb4GeTwSjXxYWKevQXCjasNU4dWoOXyP
enQmScU2Qk5EpSXljjeAIUxJ08bY0FmOHefNy41eT1FSbP2pBstc+TQHZeKY
fnLu5eRjXk07oXlyOJ2r/IUAUhtO3/kJiPgqD5Im4xmfCLZUsA+omr4G72RX
nK0cfUhH9c8rptSpUToLPAyY7XgbEwx2vAsCk+IJjIfGvp7G0uJGjBo3Nv63
Cs9Todl2f5pE4zYW+7TyMUbjIwwbIEKL505u1wQduEL0SSwxEPEV060Bk5dh
znxalekuHQ6cpDjXKk2VXduNYXLVfPxM5sR2VKYHs9IIuRBRVWYhdbaHwXo/
N3osjSBitU2VKXHBK/WBpy5XSZwv9+ksuVpcCI26kvcqx3zjkXq2DubBPhgS
UjqyE3qpXteZgAffoIc05AZAMtzB432O+6h9SiMXVg8+nyykbJv80PmdUrXM
7QRBwS/MdhswlewTO+j5xE6HCmDGI8/V+S0i8v2HQ5ZTWOPJCsizkQKzqf/V
CYDaslJCcc9NmZp5n44e8i8jlxkOi/PrfNnBlygntfUBZFGyzNPfRv5ORdgQ
2Oe+pDKW0M2dq4G9C6eLKh8mjrqgJAXwdD0vuLuAUdnJaNd52xfEzbKVUx3f
teGhVBXFluc4z6LXMk8NE1S9990JVscZ8kmB3L9G4ysjiD6Fa9F6lsHZ4C7I
3rqJ29fkvXdsmCviSY+IfJ83bDm7LuRH9ikrDVJppmkWPH1gkSr7YwK7urVV
FZJpNN2XzsdmmLWlMuG4hdz7q30ZiZ2XKBwjSZ3uWva5mB5nNlL0aJku59Tf
Lr65cfJz4BuWuD3b7U4VJLelGCK8aP+aHtzqeAYSV9Fa6LOuPLEcNODBS44P
mADHDbJIQ9WhFHLBJEW3H96onzVWrPbEIuMIXuFgCHrmSVF7hsCxjfhhz+zT
AS5Y5tCIBPXyaOn5f4lcwokIJ1FSidPP433VPnvcZS79Sdo5Ymk2XywCG1Ib
NkPle35gKPW5+6c0MmXOUc64mFdbGWIWrFV42fpG47UoLiN21W4qnAb6f8Pf
o3KWnmjbcv+0e9W8oeSTLVpB6ff2fzWTNWM8UUWe330rNwgAgakSc3/E1q7O
54eeVAJ3pqx3EZTyeDOi3wvIQznK1owKO2+EH/Ml2TD0xlruwXgUjLOGui2G
vMHfWqW3XBPHBY8VNVb4C0Ri2/+OopU3yQRYJuyCAP4j+RnSalSCp1Oru8to
c1Co+V/w7JHmk/XbpuVNT/dJMa0S7qVtreT9bVlK7VDJvgoMbct7f4QUUna+
ARLDuaCSeuRLQUF5jSj1vJKhJVvTHyatWAysW+o4SOrtr37hGGPK8bpEmAxv
wNW9wTWp2nxTQHlk8BDu+7LrnM1bGBmj4UALhQ0DoGeJyyaA7ipYOCY4k19h
3SXpBsGNjA3oQAOb1O3ukZhQHcSvRmLzzwqAIz9klEiuZypfsCZEaXQR0N5Q
mnhefuzRJwDrjwHwxEecIZo95ObVlpCPPIJWJowCMTKN77D7Wc31djHCv3vO
M7i4k9U6/ZiX200+jaenSDogGmnId2dAFTKBPRGvQHEsnC+VzWbbTQhLoGvx
kUGC/qkgbEwvBipWRhaLi9t9RrmxwfE4/9I7+2sP0sokZmLqYMB2w5ngxIoS
RLb0w7Dmw8Yv1GPHk2keT/DTpM/PTlyaD08heZcSgNTrYFmP0d2DTyyc/tig
Prn+ZkerN1wEOIJkSuI0ZWyCon7BSOmVibY+DDZRgU9Cpo8lWIR8HcQKyT6h
cX2N+Uw4mfHyixzttlPfeL+IE3xJMQ33jSXm6zaq/VoxvSAHrCWhqV12enUf
Kn5+Y47fbucL0MC+hfL76zR3zQWIbBv1yFQdyVHnWQ++HayUDXD9R3XxBH0T
8yVQb33ACgDsPhq8HH1M9s2kb1wTRpphxJsvaMo1znYl9rEX7227oQz4jL7L
+ZEPKFqDYLzOG/HEd4ptOUi5tEXSGqRJK+CBRdLybb+tmiMD44A0VCNDzMo8
xfn2SLYbJyj91+Jp2ZbGmg2HownMJ46JlUeQtq74BQb6IulkDjQOSKJvtIrR
46NTlGm6lbJ0p2dGTwRKmvogEBzwmjnqkl0vFO4wb6B2J0vUDvM2kQDyAorb
C48PNGvm1qBuNjFJY6Wd3i154SN5cS+Aik/W/YBrcHuZ3kjoBstGso9DJ6pF
xLkArm76UEHa/nqCpptEYF6/CnwSxKsEH/IKsymgJgYGRiWsZj95Ba/TVmFI
iQNpe6TMOXpHVYddIzcT3dWp6lECKIBsTN0GtQvrmHGwmxbQ0wvvdh+k/0cf
wfkbweiqb9svRRy9OEkzW20jXOXPoIxFrPiCLI3ns66de4frKVw00RitOV6S
r6T1jG9i4kc/2jhinrjGMQDZh19ri5XIZEgvc5hRQr8Sa7rCEoEXGe1lEjmI
rTVeuEZ3VPd4muaLOez+ZbUeZOWUuKWOqbf8ZDNMUVlWjPeQ1KEBWxsVCSnp
lbNvL9kSfboB4zs5aJaTAcq+ikpnDTKgIWSFTBFT5aP2lmKV67ZMv+VjWSn3
kn53UtTI+hEkplY29WRkt7GFofQJN7bZ/1UjTS64/llXwdoM8P6QKS5kbw2h
xviK3+x55m0Nly0JZ8dRzKX8SBiEQP4qQiCUIou5hwnWHxTNbKxxZ8sN4n79
Gak+UfCDKvk/r+DSrB8ioqMJ5XAwoCDgxw+LJ9D+yHjyTL07XtkR7i5rSHAO
0HKnkrEOpNz7jvET8kmNnaudjYOVct5W3ayi/2K4yVinTLbJuweQiUwff7ft
+M0gsuQwBBovnK7v/ZkfQE0GNuWSghmC7m0k19ElhLLTuhvwMLI4Lv6qNJ3o
7SHu0aW/1pvZUlEOe/2FTOoQiJ9muP1hqIdo/GEht8db3EOqnzZD41Fp9Q1h
jVlgiL7CzXRdJNxJYdqqHE5jcqs9gLRqxnOt+NNsBc26Dr9XklOtvPubWnX5
DlGPT+M12wWu45jvIxlZDrY3mrlMcCWOFIigk51HYpl+6kAGvVZ5wq6pV1Mp
EPGC62AtjM1QJ9Zd6azSGX30aypSUH3xBXHxYqoqS9liQ06ydPNGm9cOw5Cx
77ZystwCZXfEWg4XaFEAz28CZiMI6b/jw6riXNZS9XfpreLodN1KLxErLH1d
FThIBZbpVBa8lhaIwBPYLsGrjHYQfIYiIEsrCJ8hSLY16Y+4x39HVOWcb3I9
XjoeGD73iJKIC1fzu6bCWoxt5DDWeZfX6AWpwbWLW0C+lllj5At7gOTj4jRe
QKlgxW5Hx0E+t59UeHQ5xreRAUs2F1VtgI7CVqo54QoYBt5vlkFQkGnL1toh
/8dwGNXBbdcsl/6Do7LyLENxwr6cyo2skI4MeVhsJeKTlUYgHF09AvBuwDAy
CQRV0OQ8oHJpqtz8qxukBGpLabuVPPqJpy94ALeLg9UhhEMEjn5/Uaq19BtO
55Nkw03wM6skRR/O/lWYrVYj/4ZO9cnJbH+C4K6yqyCFHJatyHUdvriqZadc
U2o2tAmP9R84c6ht15r8fdEoBKLIQdhXLHgrWijYlRFE6vZ5mFYWPy41WyNv
gwHEv+nLiIFmVPTzVbkExgAYHPgiXLFnkv63CvMndP9pd8Q/KoJ8NMdIKjjd
h4Xpr3bGhm1xwG2MvIeXvfsLiGJdqqLJ0eQ/QGuCUoBMR0j7DhxQnLVJK3ge
UGjY/28bUJ8jnHJycGf68lIolOsKK0pS+wJ4xWJ/qlTzH/K7iazvRgsq8klu
m2CNYD2LVrdymzskDm6BTM7QuYN+irCEN7vue5Pte50++0LBIqcM39xTzabm
FZyP/7ZDsbNRudSpGkYl8v7Cu4FzAMgIF2YIoB2+Psq7/3gyDDmSnV70nW+Z
namWgOl6Ep9wAsP5IKjhOwEvQwkLxy4AP3YVxhmgLp78F471TW1TqKoxid38
LdBVmnBs9SQkI/tEak67FOzEy4vssHzL0VYHK/5Ve7ezz3SH7Ct+LHe1H5t8
jJb+FgOifYKW4dhri4IBXa+S7pMoESs80ZvCK4wnNH2Ov7ie21nig+xQHrLB
IKPRtJJwBbdWWh6l+NzE9hFkHpQaCvq6WcP3k8By5hPNNEiXA0M+3PKK3kbG
NGz5KsK39PXtpp7cmLdWGRapWoEZ2WJcqZVn2w4RS4/Fdu/6CDxlTAxCwMe5
NEhx+mRRiHkheECtM0nNPzE9TGFR/ZgeLp5Qsxc8dy7wLGGbMnM9mCEXtCFw
1Duks8Iqqe99UOtNRNPN7ZNhdr1peUT1TOhpUnMwzXh6fIrJBc/InmVsbX2O
5ZYjCWh+lyjTyzeot2voZZ+OzufZFhjbPz1R8XJPXztQnhp6E6bAoZ9CXCT0
p3UXrhtVeqSGd2qrSvfAaYKD2+GX3Tw/qSmKXpU1kqwuRMmlnsB+4xnAVG96
ppQJNIbWRLps3US5QMa407KiKwfxNkAqR295KQVlnp3OZjcKP2snGnNXzbPm
QMUh/rb4uk0iSKIocvWhL5gHr0+YWd+bRkhmOxKub9XFWVn9wprMNfR+DR0J
RwZiQOn0tjcRFRMvek6cGDp8ZctCpjvzoj6FxzOrUbYlGVT8eqjT8Q4LmihS
UL2YEVWyTXc2Ql9Z079+QZQUXbqKqDe0Xo6gAQPk0Nv7PhVkvmIKpkYuaO5s
f7siaKr1sLG5YkH9Wk+Z/cbWisllESya2LYc9NagugaeozTMAWLBmTVW5dbj
BjoORw8c25d8O7JgLDze55z2742nesyPDjd1zcyM3+cLiChTkFSjN5hmY2Pz
d75vpr4cb565gNCJ6v7/g2p7QVmRIJ5Ox1YCu4GwWUj/QGhx/Ow60WoCB1bY
HSMZeSitjrISmtbPgJuw7GBczW9qnbUrNpEfzrYP+jWlYhYe2j3Rf/qC95UR
F/XsBhFyJFC712ky4O89kBh74b7VF7UOFaaHRWSUSKwt9bjl1JalpXEsqen7
PtkTBiuG922hlXnwzCAB5QEMCtabzNtSA4gwl3w4rAILpPvMAsrqH2N8qf1y
okY72UoQG/anuDheK5jG9fBUd99B6fpJXoqp4BR/IvJ6hrz75PCMug67TzVh
n3YcATSCguLEGBmF/f5eJJ74W8vY3vSksL3sDJaj0XT8bHgK55FihEmtFgIT
T40gSqsLzS10Rm0ujb3BSiYEHsOXvDZIXAFgUWSFw6XTUm3tgY3GMOurKtpn
7NIy8Kxe/gXkE/eVII/h/AKL0vdviSFsgsqa4Yo6XtuF0XsXVMzsA0yoNF9N
5OT9f2NjU4hnXS+NcChyZiMoQP9+1Y/aJqfVS3h8eUi9FrI0qjPgiC4REXDS
Ctx+cuRbkrRwuNf6pa4oSJ2Yd7wg6mIgoOYvrwBe5WABV7Uq1rtn7TVvyVjF
njNO83NKNc4T1CSl2/s4Z0Oyok7gb3iScNpmIPGKRdJWsdnzYN3sqZxpDj2l
nS5haf/bi/l0hIV2qPhZIdlYgEwWMvDjZVUvq+82P80LIbsxeX76uqym6lWf
xTsyNTwvfUVFaYr/tO+tLCMQBmaeTp3YuVZ45KxsnoiMLR7dsMsuJ1LqThpR
iKKjK4wQWagzoIg5KuKLM4Bqst/XvzCaVSX0kbXEH79/r1/alyy+eEDo8hzd
wlS5UcWUcGmtqBw3BRGnJ/S9YfkbQ2eDO9GLelczwxfyXIebrZ52Imzj2J97
CdoSQTCIggMIo5rsj5TRboC4atCbLlxmI+mop1x7DfiKxV3pGVYmNjv2rYgN
IvRQkPVHjyQs1S7OIZOgtb04LR+RqxClN2XS+OH0TrzuMl7NHBDTcy+8WybB
smufBsjsf0cMUMRnHI80hoaGYcb/rIU8uuuTgm3NOTjTRLemV///zeWQEvpI
jV4wLGpt22zn2fG9c1MHd39x8qmCEbEk1AJJCDCEdUtqrMje2ZY8+ha31hlX
52fK66mSY0K1bTOJsq1RI3fdVROuFDNcOo2wIJ4j1uKo6zIp206pUV9rKgu1
G4WNnYMAJOcuQtQDHSlpMmtn/e4tGZ0cbwFNI5nSlbptByMM6BpPjmsgsJDB
HczcT+RSZVQ4jbRAomK1JmSyN3xsZJPcnLgz1+BjhYNrNouffo1d0o/m9pfp
lAXoul3pBtVzu1o57t3noKNqkV099HPnLKP5Wod+Bdh7iZWOFNXuB31/Aknr
FhhzBqHVNb1hcA45z8URElGq1IDn60FmCVDhejID7o1IJQ+RXnL89ZwJsJO8
0/5cfPklcUMMRWrYRDMNzb9ApfmjVZsPW2FLrFusYAYN1fqYwFYnRdZ7YJp/
79Y+hfxITbpxxeH2w5e1X7i2bQ5aEm9RRDfRqgK2PLVnBRJNwNJZLEdlIfQL
oXgXXPVwuWS2NlTbej6MAbrCZVrRj/tE6Akj+xUKeKp2c9ohYtwKRfraP3Vo
S/YeEXDLeWfLjIudbxJDxM1VVtDa6MMf8/XfVYHGo0ag0sjGpv8j3a8Cx6UG
U5kAfIjKuxpZ32vfAzzhjfEtHi7HRyFJ0q/r83nlqTqCzSxHUaQF5WgD4qvC
ysGjOgbHiU1TMUCKVFb52XjdKk3JKSe9TzG099zonKG4V5Gyturtfhn26qNY
KQQhMkorZLnBzjHhFs6tAPiLiz+U19hqRQa1f+/7cN000L2T0JOE+sfztRhw
3yx8l83UQsSuYmLUZTyfQW8sUxHWLss759Z6legNG/KIypnCTtH6ESj4JJ+1
GrIg52QXxdDfVFfWilqS16rd9eEZI+b4ba9l7L7k7pk203u9+vWaIfz7i1gX
6aR73ktO3C3/BuQvxhGbXTnTr+8XZ6g6fxIdU2lOKcqJYFh6PsLJ+vcyH4OZ
UFzeI6T+FtxhHuTAu6HdyrS2IYvbSLTbxMFOlKyCb2Zhg/2pzueEEBtwJg5K
rQd3mV3MA1BEU8WmPlitUYL2glF91tP4eogev9ieEwUCWLeaF6s3L2Agom97
Hr0IMl9dkynODNqZdcQcwa8vR135n8yVjlL90JsSX/6jjUdgDzpYqjzTuUXe
+1J3r00bdASALpmVytJ0rGKanmCp+nrNulG1YD5fHUMIKFL9sEXJVx83rthd
m4klOaeWG95xEq4XEOn947ThoAc5F2O+y7jl3AMtfENmJA1ZsR2hTbukqp+a
OVBqWryevVB5pjorWg2mkZHaoXiVyu5761wOvLwSDOH+cxv1NV8qQDKo0Wh9
/H6wQF+OhM9wQIE1pGXdJahjE7frhnDJ3SY3sAdcJAibw0WXixiX2klXsqIl
8yxQGQxiEvNsZnD4dcv4jbs7q0Qv7XcewLQXhLIVh0rSL+IOw4dk2yJbRop2
WLkEWiYLYbp1+M4Xr92GNtiYtE6OMPqzOJF/FqJXZP5Asevt+wtsVhT5DJgZ
0frgLbC094lP8cv7At3woI9GomuY6eQubfctIS5ecRK9AHYJc105r6rVnHV9
71vdfOd+JMuCqf+0I5CdM74L/Z8LWP2kwBBDq/VccC6rK8WzHKSMOHLipr77
ez0UM72B1NoP7fbDTL6gAId+Fcv46qUJzL5cveewfKLGMaxYrZKPyz+aRhfi
6159vBWMlxAohseh3FanY3iEwD4DXFEso8O/TRN3+Zl49ueMI3MoDGbjK1wh
RGWPRHBhgYCXiyuVsQYbDiIb0O04VHnZt40v2JNwhr2rsbyNsnzIRE40Cv4+
nCbSq7BRzvVJG0FP1mAd/fJR7wrRuXIf4kx2LYD5UMnCIQ7Fo+7PiRuQsy02
1GojkKqnMYjI9jcwxMZx7MYkuDH0QCAZGVYSuCCkOV2Uc7PS5OjaNbbIkSOG
Vwj6U8Beij9RnvJLUIkqW96Niw4cgBzPdY9PEYUrS/2WJ46o5X7VuyESsEsf
y48rq1Gbl8GCDwCgFBlHbYi5Yi2joQMtOyVe/MI5Yy/fEx8xrhAk9tf8GMk5
3ARaaOmoxpZMqyBhmWxQXuINOy/xuKIJGqMGlUppkIKr2ior4nhLfUynB3PA
GZQWBddtQCda1AfRjJPAM6obJO621TB8uSthXA2mV3ASwer8/UkGrc29cuHd
i/bir/7ysZPWO3of84CEKh8bb3GyBZRXKxocKDH8w9yows/Rd7pfrAGPGaMt
5gEc6gx3VhecbpecVuesSMS41fDQsd9pXaY8uHc/6gFJG+umbZhes4ePwTRd
c2UMgXa9BYODZVteY9pzyciuxnXsua6nE5eRjadrrYZJxpT+pPcOgkPIzUTg
bP5PshNS/Xg8gpTueznEl2QuB9sqh2yY/Wdox3i5Wg58cHsF2QgQtHbx2jzo
7dAPY0PGJeoo3xF8bDMHCzt4qp4YVOBNoqiMn5muHTgyff1T7rkrxNfW7ev0
QygmgXYQOQ/z9QtISfny9r4EC+62Dt/PnWIQ01fYA4OjI11d11/EXghPHiMw
/FE3q2iiGq1hpjQhJgntcOFeprEEDcdxMorb3XiqFaMFLpwNqnB3nVLFmHC2
bkygOfd639V0hzn85PKERwVnp4PZ4iVSI0uqxq2t9lBbQKj+I9Y7wwgAZBzE
YIcNwLD0tbUUuiBDdDP8Xvjcco4sOmZvuDJeNyAPJAHUaLRwQV6JcNKafEpy
ltyQTotSxrw5rDKhZwVM/iGvdqWtFf8L5tbRl8c3MFwkNQZYSSsvc/bWQL/L
5Z/hx4BWfFvybCnYBKzXY30wFKcsDARkuCIrbRwFOFTCcU7SkRq+yTmes1Yi
BTh4wPJq1ZJZ5IYbwGXM/3pMdkdbF/YWtxqhS1EqWi2ze+Yn187yti/xqewX
iVhZBLHhwwaqW7YpTrG07BtpkYoPZ9GCQQhEpRtD+rzz8RvRgnP3BtBRr8ph
LxuUcdl+RszA0JXpB5NEfXTFgupS2n5FfXfDGQ6gIv8OsvMpasm3jgGZTnC7
+iCcTiGwS1DNApRkxKgsveAduIIj/04FaZkQS+7LQ3xe6DV70b/NtvHElDXB
w0o/+XTnqktDbWxpkmjCnySxqzxiw7WJhXe7Z+R8lFI5LnrCKy9BngnsKruw
A2xbWFFRsCpCjvWdzPz4Fp0DU4Xam9HhvdTQ382mQedUlWrRtJII8DfCz3r0
gS9reA+OqblDQDQ/GUC5iHh/CJdEni8Wjg3CHJmkBYeoJQUHJRtTgo7lATEQ
+NAkDTbf7cfx9/VPHhZpphiKbPC6AiKuUSK/5+LG0G/DeGorFaJSOppE+YNu
gi2ZZnbWikd9xF/M+BkDv6osPe+fCR3+0TWpARQOtx2Jc/XfZ32T7pfmP8yF
9W/PdTiKidRaPaw11p15zXW9saGOcMJHH1ZYGMrtaRNDYnm5GxmAqd0uAqd/
q+vN9CoLG+gWTbGl4lIifFvradZuVQQjYD1dtVYbX8b57W3wi+yAJFFDxa8S
ZbhN8KQ4C6LT05hOwr4DPr/HA1pNrwweZB8I7ROedBPyR/CHuZDXVP9Hrqia
8RZWe/DNs9NjOB1vAJoDkCzK5Zokie2JsNJgREllU/YYNpbzrExTP+MezzDZ
utmeuZEu+Zadb2cD9dRWvY2ERPGIBxWfxP361yEU/7k2f+n0YxEXth5+S1zP
H3t5LKncwqijbIAa5U0Fgqsnhui5HyGXD3z+T4hOjXzgbkZAmBlU+QIyRa46
w/U8K+igAr5SW2Cjv3ANZTCeV4Vkm68zjImbLxgHJYytj2aanvPRBm5sUlsd
DS2YYdJgGlOZkSXD6Q++8XXIfqO8FPA5tDNsnVGbN5z3EbTphbx02Ihak7Ry
0F7y71jETnJhrt0IZdbH51fb9gggAkqv/vwnNa+2rW8JhIcJu5ZHSlAzpQqO
/m+k4bY0wwAWvwCpCsj40KCTn1oCDBA1Vbc6qsGYu3EP6VyUr+spSK8pJRke
gzc1znkb3sC9eUvZfOoFZJldwbyes2IMBsp90u3KmKxbLjU6TOzdm3KFvrLm
MZPq1FL4TNm+Z9dwV1kAGY6FDFRejvrB3dylsmIwiOCYozlM4HpgI+PO7X7X
n4T5b/0rhiUEskhuIyHWTAOSWCEniq8SbrI2rxBLD4+xAq6BpPTfJgP3GqL0
rkxImlfqBRw1F9tc1mSHNw2AdEEJTFJZ7MRp3lPEPVwCyusr+kxsOwfIBfHC
o47b/zeWbHtJh7CbyNaHl0EKeH9caaoCB77TZfKcakaaeyeBuVlLVn3ARy+2
XgoOZUPkD1xcp6i8b+YD9IegHi5BrT0/Y95+h2DLIGIKsDy7kP9hpFobkGsu
R9j2Ij+coLrS0IoKPUR3n/bEmc41ERRARQ1Lxzwu9NbBoKZhbKqLHAmuCgSk
GGTrLFc4njsDuKmdpfoRU8a6uQkSueCtWfCj8xbPAcceJQLrY57iNMoCH0sm
J/7Lo7D8RMpCP3RASym6+t3JddR2492Dnbe+tlAjwtrAfj4gZ/O3ZMcD0UpN
54+PBtNPKGo2Rhj8sOPZscIK41oNZWX9zwi1CnrJ4oAbKm1Pqj8vX6WuXPzJ
KDK8/6557BKpVZwuxcZWk/41I/CIi6122xbH1e6q9qjp3jb8dMEQCStOQFZw
GU6/ZrA2HlGxyfJ8wnTidV7+XC2cE9sBB4GPjWa8rT98LgqxnUN0px/ONaVB
n7Wb6Quy8ABTDAr6UNCr9KHPzEAkLJnrkNF7sfGRBlErNAr9EaIAoATZmkh1
5uM9PptjUxDjZMYnbTbFS7+0LNtyee9ARwue0ezKApDU4TxrvfOUnIMmjKHx
v5gbDR9NIWXix1WRBIFrBmo67LUXHC+Hit/R/YrFCBhM+VJV1x37xKZmadZW
Vsgitexwk4qvQbazTnlO73X0mEgYnSefLe6Vc6TM6EX5EeejettpzQWLbKVn
1hbxnjSKQ9SE95r0iywJLNwqEZaC09ffjPZV6AshR7pQnM1qJeGTQhuz+CG2
1GY0vgfXzLqwb26d//d83VDK8K1F2Nvz/obOpEnGCEfMp1BrC6Ro2ftwdQC0
7km390Mqe/yBBecyD32l5Qsw4J7zCZfzB5M9rUbVxzZ3qt7YCctmbLSV7XS9
3abT7s7RV8LH/qELgXHQEGIsvoZ9uW852uEqQZ23x40r+ewm1H2bzrabsPTk
rvarLvrisIe1+kWuFCZ6aPerhvCGizbrPf6pVdhp7gGCvVlc3CMkHQkcznPO
2reOWQ9JZ7MapZPg8MSaVjriZhXpcXwKHbp28p+doFHU+D0yiRXK9ImYcDI4
gNpsZH6jwZXfaPlzl8ZshUIaM2S02I8VUZnY18LK5J53TWP0CfcF5HL7vh4x
o2TyVOac/KgH3aV6S+4yFW0ufhjYXTd3n46/aQgZfss0M9kiLQiUuB2PQ8jH
C+nJIO6lrjMUFsNz4x+JTnbAqi6+J89nRkQ57eYDL8y6A/b5almsb6W2bl+G
VoRQsfM11baj2Gj5P9wO6+eNNnqEPxp/xFYDChcRpCOFBcudrDFFs8qHl4wf
VyJU1w1HP4tnlWIkrPcyPDPbwznxHfIjSYQIduSFpVJMvPcX26I9oTSA7Ulj
YoHcCm76djcqumr1qmadurYwcprVSZLvfVqni4yLpoET0vI8M2YwyCkR2rsM
z3jjqzihxcjNsflBP0v758fgmYULjdJsvvhO7PZTFiotFFQbh5dehB76cSSV
ENBnTIb67O7TPLTbK6f1FSH/RwlNif4GlqxPnbUgCUoTGOHbqnjG0YGbUL50
3hcAzhloZ++ZiYrHzaEYNjfZ2vEsb2eegaVy43w+ZR+kKSRGvRu1RF2PLXXo
nL6UtN+P2uGolNG5OycJHbKJF3puH2q3GSimZRH/OJC79w+AvhFmzL+aaDSV
tb/Yj6U6WkLT0LfuW9pjhk31nbxSJxUxA8DeWZVwcSu3uVROWtTxoKs6fH6D
WUBxvKFnlmprg33obfnuRGGE2J8l+8XpajrUkFQ68DwXt5fx2S8LIP+XLCul
mFrzZ7/gNZVgn5lvOQ2HxRtt5LPOkuG2RVGzfmNxB6xu/Nfa90dtf1S6b1pD
JLTR09atfP4knVlPEoh4zuDrrTbjRuC7N3pkXaFj+nj1kh8hVG/ccU02HQb9
RtgfKVxULCBaac0RNuikSfpzQBdvsEIxoAVLWGHEIwS7Z6NB8Mi/+iZsToX3
UqjgLuZ7rWiJ2mtQq2nYWiRW40hF5Z8Xyzc22pDd5lDI0IQuO9YuMPuUiz6K
YIca8d5SXU1XpaIg20Red+UCF2sdsiUdcxMdrIot9GF76WZnxc1AgK7cI1F/
JdOEU9ZKPqaXWZHNPGt1daQLJAbvSlELc9g2FGmLx03cgdrcBKUuoLQq7IiJ
iDpTqvD/zWRMH8pIb9eANbUrKgbD0IgpArypOUQGkYn5vvt0Q7XX+lc35cQD
2IdBIo51ZD2aMb8PwlJX2kFHGDu0PBN9zRAyTPeUbeiMA7pMji8SmcqyE79F
qPiWGTpxOZaFmPaJ3OzYBkXdCU5glIVLkpRy8J1NrbS31vLK6yiVvf5HJZrE
6qmDRTOjs/ibGOa4tEEF2MqzOSzEKZ2oMpSkK+oU9NgsQ24Z3T1wRyklZhlv
NJHSfvMlLLZrZOmiiIRR4ydRKQLy2NrMQiq+XTt2+m/wSLV2mFiUFFvXX7lc
Q5N+Iq34wBSYNPJ2oCX+gB5g1SsAPNHQZvFoqxOfEELvsGSo2bJ9NlenN8H5
+iqUimY94bduyXVZAvqWyhnlr9/gkG6LEcAN7WhUh5vDtqCEtKEnyVQYrVM3
z475c2lc5lRolQbWEH33MKPLBKCHvnakSljWeDRGoNAbmE1ZQfr5R4pSOZry
AblqaBoFgnUqtyI1W0QDBrFi/LHjOJa6NOOAuJjH019JWtwf0gfr5dTcCltN
xh/k/AHAWuB5YnkctN2UVkp340HsvP9vNkycLmTRjFvoTSok6nxzwLOnmlwC
bNIKYIqLDSmHcNbyLkA2tpck/HUINz3NT8CoMhJt+o5V5d6mraqr/9vYj1Pj
tbcqm+06dNkqIzvoURU5qjb2wxXjqDaD6qGpLwHgRqPg+yZmjnLDFjJ690G6
KyTb18eGK21ct/G6Tdx32L+Ztr2kueEtLMYmAb8cMhdIOopPvsnflNo3+PTI
AGQ1lV3bZ+rNx+ckQyd9YcttXiBlsCmFUMcVcP3p+boAGq5/2unZsp7MU4cN
zmNtBZx0BXS1h8iBdn5rrB3BxPdsr5UtrzxbPTih5FVkcVHh/7N9IWdxzJsV
JoPU7xf0j7vtLLmoLcFoy/wBZCEaWIXZNroNoHYQyPnGHEuEujMJhfkdAHJJ
/pcpL2oq3+NJwxu1pVVRj3zRSgn7izpF4HAoBDO6YIgr2aUVFhSc91urNrxP
TuU5wZzWLipsBVVgXnBQ0dBWzdFBVszxp8vkv2Qn8SlJVAMwW35Y4065rxaf
lggj+T9EzFOBapvbiuNoRadAMOFEbDBerKdcnjGlZxV8gYkxxRnDEe8Wa9Ja
ZUYL5RQvMvmnp4ncwJd4VmUwiamPER5MsRM9tfJXJ0kMF0RL4rKW7kQJ9iJe
6Oyw3gsEps33Hw5lGkGnicjXChN30ZwSewqC8WCD34/ylAkRW6aR6oNTtCnL
jO87nNRkLI7fQt+dpoBC/M2kb/UpikyKth5djt/tR8Zamx+F1GPc1aJviiKX
fldP+58F9JLImIpfYfp5nQODKC3W7xjmrjJ+0qPTElRO13spBkAH2dBJ9/Jg
r+F1WIp5+k5FXyYNmRCdTJFvLCUB/IomXo65uVGlX/eT39pL7YmwFJkpY+Xt
KyKYMmPBYIbi9KJOpdRJXJut1SjDy41PUWsfm1aFQUOIdn6Z52LauPpWWiL6
eZ/69+q3ISqGKhzR0An/RwV/Xrp8rYVnkzKANiYEiYB4SadYnBsnXXHndqKE
HIQO36oEoaVJPSVAGaCDqzdDSjM9ptjSLfwCnEp0cOt5TbhVJNXz0ToV1or+
wGbyzyku8vnftKxdGn7mGk7JOpT9S1t8MOWfewuiLjpjgIGnCd6zhDOEHebr
ay5JaDIQqIF1R0kkjJE5nd8fZ4XFEP5KF43X6QFL8AKv3pCzryGXCbc/ar13
19wl/KGRrat3wvKALzHKzKEVRSMvYGQL6ENjeueYTCNTjBD3RbKHz2DvIYU5
SJ4wMIPdE9e6pbv3nijPsK/NK66KjaaIvmepemIIjnbU4+dBaGZkmRDT1Rd7
L4PmUfABCxoi/zOx+CcPndHFSapd7EJi5UiwyVA+Qh4+dTg2V7Ddla3bA6z6
W05aLpLn3+hssiM1jlR8ZJWLy8JhoRpxLaItEpnpYA9/SPklAHpOSTpZQRqa
LY2Dqszrzst9whoLbNiOQgQobgkwCLRbHiCFtEsZwxEGnG9NvQG5LTJ2kNBz
At6tUxFVz2PmD7SQyip80EF24Y3zeA2qYM5JDaw2GbcawETbmS96XuyRq+13
cyZF/2+ALaplL4Sj98ibsbjKstbcF1dRx5Ooh76/el7BDX6U16WqOGAP2OWt
ldMtP2xsBRaMo8RCxv61q6zzqJ3LCzODXxv3aI35pTLNhNdmqf9POeLzgD6I
w5/IH7Y/q9kucfY1lg1nIcWrvmDUe6hjYYCuVS3PKWerqxyauMbXo9FyaNTB
hIo3mwpaoj8VbGdBZ2RIzTNrOmrFr85YIt9l5eli2V/kGNLs5TU9sO6heC4o
eDK9ThjBHJwhCOR20SvCWfz+s/9g/lBDIAtIoLNN/NTXT2p9EuNwxR4lznpd
vKsmasizH5FZ1iesYeSABR5X8N3KoPRc6UYFd9SneR39xLrNGsMoLSo1u3kq
7mHPgcH790W1fvkBy/hNHr4zLBOUBD51gUmgCAq60SyZeWT8dzz6kqHWgF2F
BEQWKR61OySaHe8kXyodpdWDgLpkJQQGTIvUt5YtRjb70KMRabAigeHsvI1R
fJd9UWFE7Nr+4KvKxQ/H3sqbcavT7j591Gnss9Abw5AOyeurAlH95HZFY6YT
lzzlIE1SEuf5jn/zfKArc6WQPnyQApXcAZ58QlbhGufsb22+5l+xo2i+9yxD
tayhICFZCrN7zD+9zUn1Z91UrR9fY6633E/3qGZ73PD4X7HzYpBIDIHwb5kZ
bSVdrZ7h7loJ6ZqeFbZT8mOiOmbpYJc4DoWzADFUqhVuvwo2KlxlLjNUACjk
GV+QzNfb/Bev4W5fQ8owqvj655keHGdrJIYD4it98LreES+TMHMUhbXJ/puC
syQ0ynuGJ2Z91WOn/evf6ARslztOib9mbpnRPpax0iF+88H/HKQUxcVvV8CH
7oCG9Bub5KTlZBAUDhnLMDAaf5BDM8k3vVDpB2ESTp9+fs7SJkfxn405HXzv
AJQxKt6DLcxg64Ar5JM7n8KJYcvrAVbTvoSTWfK6d6kDjArvK1VguYCSOi1J
fuYjOEVl3gb7melBAtDFRuhphruXOw7m8qS8xfMExA7CvQr5AwKx++1/Rki3
fr2iFj8y3ZHT4z9xLLa0PGoAlAc/zFAlG4wdDGVqvoCubyNC/wtVDA3kAbyu
eNO3OvLngmTGkGDHkkzguq7YQVQZyR17PQl6bNKvLJhw7Ar8IMzJ33ALuhrS
UeIcFcH5fmoXL/ri5sW2TzOOXu4VgUP7ffVuj5uiLwD1M5DW4zZx5eakyw5/
IXoi8kvfbHRsFkcYK30b5inkx+edWXdM4IBc1E5ObYbEKLgOqUp/P+841W1M
WoexDeosAHsWkjDiYRB5u5Pu//STky4QhrBV8EL1jnOTvLLYteM3qq25/QmO
z/IIUQmLbh8mzOvVjXYD9PtCiWuLH0gt8C2j2zjBidrqW/pV/eqzcqHWnKGE
+Rpp4oZ9Pd3307sDBx9oJ0e8P9vyM/sGDnoxCXnqqc1EwhYcfwWa1S5VKMFG
dvIXqXf1JP/LSbh7jmyb7qVAsQQKwIw9j64oBVEM91KkYDSiSabtZV7U7CVg
Dyt3wqryDT1UNQWO7E8f4VufAREGj+Z5TlXjLMhyVbg87Z9115aNN1GHaN7m
5cgG8KCF1pWWicZQS7ZJIH6OSmh52gbUM7tCVTvm8KAu8a16J6FTlitP33zv
xRXfUpmaOx7y1/ZipYzt/AFpR+ItNS+pAAcwKoQB/jH4E0mdAOqHnEsCfr90
aM+BYcRrBZQQ514/L7O/C44GJgIMRBruHYUHvylMjNks9Q3LKmRr0sQfYIOT
9LSFOmrHovEklP22+IScfKpVPzdQ2BRUqY6OQSJmj5ySnsLns1YV8wgXG4TS
gJZB358xrTD+5y6LG6qYIu+zEoASIlMDVHQ/vZfk5+mYnio76jCsgTsPDGje
IiMATFVpJxt2wDPL3hMtRlV7tXaIhPox7hIEGVsjaAfc6YuU6gxZxgkEWjKM
X6hi+KE/tipEp17UdLshcH+er8sbM2YQyzBp8ZiG9EuGQZwtj5n26lWn0z10
YnFVRcCliWX8k1Ujejar1RVzwmX1ej0gIFAg5eqZVvGwe0ttuKD7hsEbqKUQ
M44Jz3WqgViBd2Pc5frsPU6ys1j3ENyqYpA/VKwFXeutqkQ9uwc2uXZC9AGu
KcuNfGokNzv48GWZZDQsSsdJJCj2hyMmnul7wu06VtXieqZicBHbEp+vSzHe
JlS876FHCMtADrez69WJ+Otvgv+/kJCaFQgDHeJyEBPecMw+3AuVHXIO1xWS
z/02LaN3U9Za/L/GpOYBKeLv8X87U2DMMMyMZKK53NGXo+siz0mw3JG9D0vi
PuHLXJEAiWH3uT0+0Hgs1GsRnp4RXPT7q3hYfnJDC7xBwRZF5AkX+I0GW4TE
sAyfvs9ASwBF2JP98VdGnhMDtD+XfcwxB4ids5bFb7Z1FIO2edjcK6Wi1F9i
IzTc3UH7Z5ezxuHsE/Yz4UI2EOw228alPVpRkF1CCdg02+CDm+W+YtPRXvch
n/s0VcBrZReDH6/tEV1HHJgai9babiuz8e4gnpPnhUVIkSzUB1CUPjV73+dB
mewhYUb6LVJ+xvvHYxHz9cSQ6pSGPdxlLLpm5Nfgf1ZOFxcOEeJk3asvfXYh
iMhxxW/Ft1fB4PYayS11p5HNZ+awbaT8GcHvg/Hvv3rhwp4ecml69hgpdfLD
mTaDz0HY08Q0y7nzE9R8m+wg5C1gEr8PHl9u7wL4qlpcbWAzs0oDkKYZWzN+
Ry5TZdKM7M956dynFlS2woMrz4FjTU0q8iVsRdLMjZlhvwbChEQVpqYCm66a
eRSiH/5j0ZPcm9kJTHnTcRVRihFMsqB4v8Wv6ulxAXS9wk8NCNrtUltaf4hn
HXhRFi4MX4nuuF+8LdwIdn0rgFLQ6SzIEhaVo8ogKtGyDlvNeoUfBW4FU4ai
FsyoUwz4RcYv7pJlVmCDt3mflISV2NUeMU5xQfAM2IfmRt3of98FwyVJnepA
3RH2iX6KgwHJfETMTJCw2wu8pStTozmeYTOh47+DoXRTRUcxSh+aCXEFZszi
3TvcO2f5ffSAbkwhME69wX51IeW1Xo0cRR9LHH8HGE1WQIvghv1FPK7WngIS
54IdjiGm9EMejULWBK7TZrf/N030RPzX7iYGINbhTfmS5JqpdVFw7a4gQcxh
kcEZ17bGp2c/XEDxVMEWgRpIzMZumtqd9GVP9VnUy0X7nDkHn14Mw7JmyzxJ
8h1izEwhgTsqXZ4JwpgSk4i+9Fg6Bd24QMjIholNv8eIeZejJ5rxa80WaDbs
rl2kRcax/UsD7dt91F5NtqRX4LPXcFgFbn2CWiBt3WFtk29cHjEjDI1f5c0+
nmywIKTIN7i4QckYa+100LoYGxb84Xk3HyX82TX+FF5zmqsWlvqUNPgqPSry
Eh5k6wdCIxHvYmN6NvgqxMNdbWVIm3+WTgpWjqL+KI+C9ATxl8wS/TXwPFuK
N6SgFVH0iwqdIfoa9J2pPJah/NnX9TcHayRLVtlK2A15oGKLqZ1YK7KhUF88
ZCkiIS4h4ZN7HCJHZjVlq5GNZa2+Vyrkuk17H8rBW1tIDQOxq2if7jNse3eD
b2RNwFrJ3T3L17zfaJiAffnMArm/fiNfoV3k0j748xIDu58yVjy60o4SNffc
/NveQ0uyrSJY5WKYdK5b/bO/QVaYk0DpJg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe76zcG7ob69FfwM1XNDTmXLgBtOMFjh+BPks86JUei4worMbcjyBRYG6qhulYocecx3wHMQlkvbJDdFb84uPSqWtal+cqa6uCbFe/roIrwax4z1n80HkNx4JCY+1zSGSbYECFFnqlTIlSnVeXiuPcscEaoN4e4VdeMv+OeVqSmN/J7oVZ8qORCBggc5nnW+IUR2r1Vn3jhRp+DVqphAMAxABY/+DReYyUcOglYqitsaXOyv60AnWDlxWxeDymIqy8QtmdCZNV2Rv1hNvtSS+/KYu4HwTVAOtiiCcMd9iZs6jAAy57bDRpPPiEcqOee7Fzvw4Jygx7gHbXIzFfyJfJkuvA1xyLxseQBn6WbwXcHR4/n/61TnORli644LdWd5TS86HLO19QFXj6tWF9U58UZOqYb/6vf750uag6xRC/14+ElkmlXK3gnCnKjIhY7fuM6JYzs1Ea6XEEqE7QSmueRgqqvp+A9MLpA5WCWCNeRq6CKX78VrrDz+Ww0Tx4/b1XxAp8xkJVJHEP0Ye1yWpD2RLS8ftcLHTSNUAUmQLk+BO7elQitkg00xA0alhKrpIO13r0j3UFqnae4/YKPvfsjTNysAL2GhGpSEaOXvvu98kqdd50XKu9sI0Ed3zwqG33gXJ4c/MypflKMEaMD0k18QrRASjmAETDwy2xGoNRcmQpR07IJrFko++GuOLAaSzhvsJFDJYSKxOyDHOsfxiyqs5oXqh3k3SS+ZRy64VFz0l7q9D5ridhRylbo7Ja54NUjc4TR68gTXPVO/iBVEWJjzd"
`endif
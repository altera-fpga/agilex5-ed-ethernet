//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xhMJzUAttcAT4oGYF3gR9CE8qYQ7Tsl08K+ctEbzpCZJpiIqJcO+mvSrREAB
7y4w/lI8Pg1isFikNUJ7al6HIp9XvJwfqRl6Fu+lCfFqmNeBCKE5zPB+I+fs
KjWt768yWYIdaLuaTekqa+RilMpCwP8UIyYO+zIlcZJT6si/pGrgiYoTDLZN
dTmZiTdBbBm5O43bzJGhFCJtcFgmU2uvJMOphHyykvlSEUMtrT51Y2m5qX4z
lZ717Ud1x2q9j38yO1a4dKI8XXmGiKlJBWfmVgrJSX6umE9kOjGxZiq8M8U6
CM3q4/7w14No9LVkWxWSpBP8dnnDubKhmotzkM9f/g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H4rr8aemHrCNoIz8172c9ZH1V20HhcAkDlRHMH4YEydDEDUCoFCRQEDl6xSs
8MhvN5oYn7gZ6+hOCUj+gdBjG2VZOXtw5oypL/QzkRxGHWaLMq2Saf7QBDMA
/uD089L0LvOdK9wtGmcJyRxjSn3nu0q3PcCeTzOnzAYu/Kj8RVbHu178r/PW
r/nIxZgzHwBvpBhCeBuAreJJhD2DtxCCjnfTD46kosDP8H/HoVSg7KHWvRyP
m6s5ARr0efhxmbp9H7cCF+CLjtxFjI1C40c/k/iu4Oetyrlisw/ZZV6GzvxX
XN9jIBezexyXnmN4k2+kJleNYG6pfe2doaqr1hrMJw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Kh00NkgxIZc0SiYjE5F/2LKK9+Qbnn6YLpwW9FA9lp5PCOZNlZEkC3gudT7Y
HrkKEa6/IhJGkBN1jtyVDw/Vng/pu79DzLFk+GdDhLJGa87oQ0eGazKsnct8
F7ILdToIzeqkpnT0DNlz646NGGj80lTyb32xrEb34B/pWzf2OycOKQ3v8J2u
OtKMGMXhVtHpcU05TvXVqEqVgf+CJCk+GAXsLZsh7iUCwZTR6LolRcfKtfQw
T8vzK1vZPGUQ+32tHLyEm6aH29y/r2y1ngIFzDwTOJ29r+XQ7okH3uorXN7r
GEDttIT1eWoHA8nPdo/dpzYo5r9oabbFT7bnCW+BIQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XZs4N5azZlN8Eovwfw7HKhM7XxKBFIHaB6YIoxF/GlF2dapp259sSz4mUmZT
Wa0VqVr2+qHOhJsdjElyN4/cidUbwl0AgxAgIuL+auHDs/oq/4ky6NmS8NNX
Q04vag4LZnFPPthOAS7R0N/TfDSGN08930ngVIkm6CPDxmyyd21uSuRpWx5F
x4Vhmf01EbXE9zXvZ8iSVUtc6Y+Q1MopS9GLIKtXCAdam+Zdrex6tU5RI+ph
H37u46ZB8m1NMOAHN6wBhFo5DXlRtkBLnp4u9RansMATIcmC6glJPrlmiSkc
YT81eldej/6h1Bwgmh/uGOvBJHum366Lj8UGuXHaPg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QCtDyo8hBXWOB2355IhwC9YjPn+eQZSUmTccLtX+m0H35QX6csBwbJ1FPnCS
mNWDV5gNRX49vXoPGL+7LgzWy5ZfCY1vxe2hOJNenK5c+fag9AJLksV6oQiO
573R5JMe3GlykrmO9NuWwetRqbDCps1nSbbwuvcTOyfKZewDkcY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mVe2W5EovVesd12Vv0rb2Lz9H1JHomr71nJknRYPbNmdZ/PjpiwUAVmFI5iy
pGKhTeICqvgIR7vkVt9pxKulz+Pg6epuzCVM/qddwzZox/w8PsHIPAnr9AMa
1G+Xmm/qOz0N8QcFjtWnnxlwzGnyZ2hL8BiBL6T4FDiXzxQ5lvCR+sJ2GTnf
hxoxklSb1E0T7I/rRnWX+u0H6JRP9vFXe3/y8XvJz7AfzJrH4ihNbiKsulCi
TB21pDXhQdPJk/TJQHA8bcUR+uF7dPiKIiw1bsN/riMIt7UlKhI7lhY0a5kN
6klZFeuoQJpDZKn+N1e+x0iE+p6wZgsaC5MrN45mgJ9HoDsAIe+iUdWng475
y/8UKmR0RQtY1NMZxsyKh9iCVIcUaRge2c5X4qgZnKkp+dpUczUaoBKG6wFe
19LC5DAVttj4fvq+LRoU9Ki1LnfTBdEQSpkv7mRKR8r67gQ13H+CbyonEAsh
d+6YTLkrHGoQ7ebQtr++WMbICWJjwwV0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eyfQe9ciqiu8Diz5WRQThUd8SWXP92LkDlTwPmA2N2mhkXyMdwwVWspeRVPG
0ubopgnmO8wua3UZ6sF4OIviCBRRfPARXWw97MiwEWIeroUgZuQThgqKUj6k
r7/PdajX/WUZ4GvO3V/m5hUz0atgGYP9qWU6faX40SUFaG5fWBY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kW8fnZEPJoV2pfsx9INAWqU26iyaQeXRqSRzXuOZE/ow+lxhQh1kRUjsWpp3
vXij8zU3JrI60AFDq1IA6LZsiav5KxtbA8NxoEljLo73enzJo3LMJcEsvIGn
7lnxnzJCvtHgObSzJq+q9AVsed2D/Ee5Unyy1KVlt5uRCqTy/h4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2496)
`pragma protect data_block
n70o1/gsRvriA669aKjqKvw14HsZxfw4y/C3B2gJZBoKOV6ixIGeJhMqkVRD
r2mJ0v+fqUr1WlARjTiQ7P/ZF9PojKwYlXoShjWH7BotOPA2y9a/r1pRCZFl
ASy3n8XaJUvMcxSPv4H4t6WivGwGhZZGlyHajJ7dX1pTSxacUHKBHdTzG2FL
1bejR/iM3TKRCh3K2IAqtNg6aqIuyzLJvHwzs56H3cVExw8ILyIU145GKKjO
F/OsWf4VDdzzc3LylGZfsnf9wRPsu6CVeVUoK2Bl/EVSYQ+WaSnDqkiE7jbp
kF3rDZ2MHKNAKPR42I0VMCbs1jC+gAkxcrzfCmlyXe5//mdU9J+TfsKOd8u8
2tybpxF6VASCxpHJIgmOD2dvJXIYF803SVbDB91TB6xMksnrLdc6fLqq1/OU
zX7/27LTywYjooxdhUvggfi8eWM8fRa5M5urFbmWlvI0SxEkeG83rsuKMmkj
tSrvou6ET91YICE7gGO+fQqKqGmiLJsdY+tQnSxzXeQNXx8HRD6QyOjwRO3F
wLD0LJBhyUGRhza3mWoh9lRTjci6imtJpPOyntIDe80AM+3x6zwkP41r3B7u
tBrcqwhT8l8KXrTu6P6WPEduso1cB1sw5uYmtV/SyLZrv+vmK3q3kOoQr9mf
b+/f6iRFzsfJpLGBBuHtIe3yNGgV5cjJbIVCgS8FPyOW9KX30dbmZ2Wt/rRj
2UQAE+f0g1gvTDlHlE8xqjUj2FBpi7HeJY+1RbYa53pSJAKmThwVAZb5wRdQ
b3KxdUaDGWgM8SLkGrBiWPuuxIjq9hvEMmSbRYam5CDxqfYgLqBWpR46vS6K
YXt0sGsb4vdp07DZwlYnbnxp1YzLLtEj7IaINDyVQvZyKRlQVQ/285/xvVat
4xapKuOOY8nhfTZDuF9IKHqWzLlEf/1F6zRveSX3ztEDGsXWtDx4nX8Ahp8O
Ho0ioaAsa+fsIpW41HvobjiIgAKCoisbAhzkZnwVNX6UHGFjxhcBjbPwbS5o
gHQ+P4GuYaoI39ykQ0whrqrIENnO2DLl1qdAlN4RsWLDpe5yArTYgTpDenYS
ZHhN8fhkS9dBpltn6Or1LmLWeqOcbb1/Uv50pI7kljIPKDcl/Fi0g1QjyuSy
MsJ92cHxFBbT2+0n0fdYsfI5umjgDoAH6OEX91aO8n9caKuXh3nituNYOGY2
kAy3qwcFRANebJVDH5sc5xjtm2Gt8RKprYg4eQyauYER0GCxqCQ4atJsE7MM
KltgW3uznL1AXUq9CCB0FpNZfb1yQg24KHIp9QqWUxAU8JZk3GktWE+qnXlS
/t1HuT8WZ6m7ey52GvI/jjfDaMPMGy4gcLi9rRoHZ/Zoec5eR90XcDfB5toZ
VOLMXsMgLlqjDhmtf65lxvi7Qi7laK2vIhjn49RjfdIqAe/vBL0i7jSyHR7t
qUNOiUCG9Fxw/jq+iKjY90wvFr1DO9wgq5pnpUKqHfmA23C2ENUfH+HmHT49
E9ZuTVsiBAHf2aT6Cp4UE3Kqr1QZlWUv5UMuK7uWRZUxv6VN4k5Y93r/dg9R
ApualjjFSyq8wdW43ECnvyd3lqly1Bz5x1gx4JzZRsvDbkqQaCtBGD87sQzn
mXGrmYGMc2wUX1yHiciZWSIw8DstqIclW6Udf1HO7g3GbE21YzKmyu7cTG+G
VGdekVF6xq3xidrJrREcpr9r+o9+zpWDt5ztgShJj81IxAc/duitFPM/7hOL
nYgFATzMzpVQjYRpLWhhxQTxbwjWqB2ylhVgmki+R169TvhGDM7qTUggFDId
ChSUWHqMKi/u9op2yqP+KGnJLr5316Sa2snW1shxwmGBG9QXG0RXztGwOT8t
XZ+sO1P+G/D9Xs9s9wALMg6qi5FHo91+X3nYYRVF59WYWigNInTycXGBq946
chI5gE46nTJz8CQ4O4QkZDZHC5E+61nWORJAYhElkRlYR1cSERF6qgJbBQoS
ACHrnWlJF0KMFAM2gpYxONu5IUjIB1+YhNIbFkEfLoXSZ+3GnLMa/2r9VYbw
V/qXVxGm7z2shLrHrbJTcv1SO6iBns+imm0Tyo+9PO8mqDi854h/I0eALeaG
fhnjM41y1I8rsgqKKFMsqDv9SzeCnZIqlXKuQFJ1hbRi6hCehhiayF4xFQPg
5r3WR/lD07BzbU4KtCOJRpdnw8Etr5OmMj29WT/R+3Mb8r6+nu95ZjCvEHQV
kIfBX26I18mabo0G1NVN6jTkLgC/N5tKJwSlKQwPeEV6s6lyUX17g5PR4zxI
sK1xa3NuFCkH8HJZ6US1Q5iTVCilFMfBihc7rhNx9s2FO+ulUfrf5J0H1pVw
yYOj5IjigqHBI/TWxm+AnsPygYuCqJPgKOjEnQaxnOnUBKhO+eeJz4ZLLinM
iP9iMxxGA2kK90W0+IO4cE16lUOX0gcUVhF/tWE0uA3M0AIBBJzj+IqolI57
Ylk8KsT8HnGeJ2uG0qSsZ/bhLHq8/Xxu7wPtDp6TwEJdseohf8vgq3GQjGYU
4pqP1Cmz/Pfz22LuLRGVz4snUdI57Q2KrYsCh25Bk+cd3cb6RE7L0cK8S7Tz
/sWbzd9zCv/f9hXuCOczGCx+QXeTrKr8ajC8a8qNFRSjhgM6a/g8I+x2uj78
ls3mBaokbkYV72tkSwHWmgDiFBSJQbmOnujVtBENLkCrsYiJRWSeRv6wQkC7
yowd6mza7duTGwBfuHvw5MkpplXYAzGA3oRIZhkMpK/n5HXeFLIQ5mkFDuuY
A7cpPPaqsYLzj/o7cbdDcwF3OQCeuG5e3BKf0ZqpCqz9G619gTxNan3/fhzW
0YQkMEzTw9pPWyIQaDTcDtU+DynIg03aC9zCz7lC53nD3C1+4WjqnvnW42ru
ZX5cDAirUON9Ur0Eg8pI9sOvjB5qHx/9Jer1ZkGkFXi9CEPPZVRERlK31sH9
xVsdjhPCHx9d9jFYtohLv6RUzme9ZcO2m3OEEYgH3eELoy9cpyzMIRpwtvHa
wWu2ohXv2ItAL/MDMNIrS/W4Imxk9xwJvnAcs3p1QHyyucF1A8u14oNwM0oM
D5bys7kRwt+LxpFa1Wfdz24qOMfoYZpPljbT1SNlgIT1j+CB6A3SA2dzgSKX
xoEMXNxTdUil2CrvI97PcTgbmuK/z36X1Z214VCoboODoyf2RPuTS6ybhyab
i4nDom/vVDaXicmzjH14gVh4zbO3HUuKoBLZmfWZCtENqcGaYNsECr7TEYnn
+HpeD9cmzD+ysPvxL1bMTyvIzxEOoOqc9KL96fODFcSzeJWJG313xLjjTEBv
4A1ml75coqprbfKH4FXKv4LFSLtW

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe74Q9QM2jdicoLC9Gbi9LjEtuu+GwDylRVQMi2UG1yYbgLdOoufQRfre3Y2dzTMyYjB/ekpdLuT6xXRELZ0YDhm7R0lOD1ujP5r/KWqCY5c70qA78s7QwiTvV//z3Q85/Tti1I1u3bioEIIVnHZkog/QOKlE41LQSL2JwYsozOOeP1pmvXR81wK0+V/v5aH7ZYg/7E/SIurepFQSkjBUdT2r0UoD4VCEG/ajJbXsMFhXjV0Cksc6leiGvYvRgrLkxt4vGgXHDO1u2SM+6WKMGvOcv8yKGchjLEdAj2e8/2hv8OVS6rM7HPae8RAlVUjCoFdd7myCXhqe7NqiOEA52kexhv56zGLlxAqYCyNqp4T2z0EJi1N5ABbE0npMO+dEPo92iBpbCbvNH1NWOg7yrdIaLivmE6s27z8Grjfc3jKoSj4Af3BafMtnqQ5qIxhFaiKvP3DFUaujR/4PQfj4vOGkYaG85DlJWm/6xL/kYCEKxEMiE0Aq2zgaeTExyrbEWrraHP3xrb51FfUq84sgZriwSOzs/hhRFuCtNymRb31/XeRckZYXblJQQ+Jw3nbDT0/wkkdG2e4PelzdEMm/PEbwN2KG+KFbIvkf5Ml79e6wFZ5B2D6ZgJ8CnuS0uImQXQGRwg1MUnmtYxEZEdVTS7wc2o58EgEyn+uIxNp1tBpNyytdtFBiKIhR3niL4N63Uhm2g/iJvZHc7Il3sZO+fJI6xvSiWPXJnOO0MmaYGCRfJwIKxzTMijfEdbbbO+Di7xvoL4WPw8PmJ1y6nuuMhkX5"
`endif
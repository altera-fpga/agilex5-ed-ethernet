//########################################################################
//# Copyright (C) 2025 Altera Corporation.
//# SPDX-License-Identifier: MIT
//#########################################################################

`include "sm_eth_virtual_seq_list.sv"
`include "sm_eth_sfp_seq_list.sv"
`include "sm_eth_base_test.sv"

//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pAaHaelOiKJFLwTPXknO12EL+CVWCwambjJQMtT5Lg7Poe/m3n19UtsPEjMB
CyMJNmrGXajxURwqTeLgizC1ljcFVxTVxcuc0Nqo5F6IFsS505uagMZedCK5
+gr402aJFHn0gIvBLxXkSvAgE5Z/jB0uyyK8yU4aG0hrsdmSfsthDUBqZJYM
JqRN9M+jMWKqCcIJ2cCvFDLfUtPTzn+ApPTF8VAygcr5TVHS5rxCOWrSREzN
57mIDbOthcnQQgHSq5CJhfRTnaEmgMB+1qQ8a9Uy7UaxUhW4sIUfbZUDWVuA
UG5iy2MNhW3iWDh97YbxaFV/3uioOkQwBiSFbvdgrg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OevzaTRiy/ywl0mrEQV/cLMUeznF0Tl75QmBupRkuyn3Rxu6l2Ogdk2W9Ln9
egoQV6Fq8Q1rJK/OBrJUd3n4ivY5qQR1f6I8+aVDhInZ3acpVDFBc7isfBjY
6JRJz4vrAWjdcD8FooygQ7zCueF/Beif4/auvsgpgF15DF6bs/UklBjorQAu
RJltaTd8jO9zOPsbZqQv6U0JFZl1Sse0Qh71OWURJeXUZMj91zdAfyf3niCt
yEruRd2Djrx7KOogmDa2jqynHmxhDNr3JH2wNuBGdk2YDXLAJe01daLH5j+W
ajxdmQRiTpM5EqSZBJl6Jg91ajbUywo2P/drlnwwcw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TLaFqWrG8cZDquievQV5QW+wBlh7vOQJk6NUfWMNoZ23GjQhSLh24RbdgLha
HfZmwFg/fkfojB8Vx5CpoJQSwdoqIKz0P72Kt8YdAsRw4/tIe7K8Db3U4ElP
VWuIeLauuhXvwCFEAW1Nq6344n12Lnn8lj7R0gnAwRz+7D7Cjogx9OpdncI3
PgO8VgfHj9QCU/8WeImmoDXS7cEgbxGxHF71QdnFUsZeLWpjEaxphGPC17p3
LzJmYI2QsAvEgATltCejluad1kVt2iYYIyxpvHlIbVe7vzWuOXgO8mOIFjEe
AW6AA0FhmP96vo6FfIEeTuwDd/GcgYQDPWlswwUTbQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kLYBUs8EQ2JHfeYYCrKNRYl2feij7eYs79EubO+djaO06+/goZGh/umQXzjW
Is1dTtoXoJgAs4pkIBDPb2KZPOPON2UOn81eLgcUQh3klUpK5uhOmvHFzvaS
Kb3aV/KbF+WonWSPt3Ud1oUAd35V3Zr/T6PV1g0YuafCke9BxhB7ewAT7vL8
pifjUPi09V8kvjktOvbO+PyTzXCc+wYh9HuRECO9HWWYuibNU2QhV/q+wpaf
1tPfMTqkyBKaOl1F07Sn/edz/JjaxY7xeT8upxXaj6f2I2ZGFqegZ5so9Llk
uM/Uc7rDJy+JtPdc+G1Ds4t9xjSiKLpEij2/toL3EA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rD+I2zesCM+N5d4uYyhIk4p0uCGgF+axwQd3VtlH4bsOSQRzADJiBBAEO0eZ
a+QWVxJBMJvUGpczf+Hh5tzemNQ1OBnW+Kd1GJV4gO9infjwihwWcvF6hKm0
FEbwLQ818sJNYS+rfBHdHqL2B3ZDBnODRKZdeGUOGzOfUqM79lg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RjGzIzL92uPn+Dtcu9umfWYYTzQy8tyQe/shC6eYMqP4N9LpJTbGMcgVR8c7
8iY+ft+FoKpy8UWTcuJpru0v8EPDs26TDdCYpfHuxfrfkOIdikCTM3rEcY24
gOnBfLSZ3lwRfCGSXIZHT+FXnbR164pnVe/Yh80BHILjClx1QNz/6iSqaZS2
mgczJPZcNrQRqIMs5Buz1u39TMnLRmhe0w7u3/bjoWxUb7rTwxOD6mUAxhzh
LYvjHjYsV9wS8aqYxoCX/ppLbqBa+UuyhstjiCmKjLuorNudZbXic3DSgvIQ
4JeEZp1uVcnFmCloe4EvMB6Cj8484NhKB1s/JjmpbFcx2OaIBgHtRALFT677
z4lVqCmphRVx5WAzFYHn9/Fl5cmUJruSbwLWLSRHhOUcS6oPYtbuiYMMMSH6
PmVBw/Rd19NqW3CPGJADHc2F2mKfVzgDgIRS4E9BRr9fcuLmqNIM7+7TAPRA
u/V+RyHVyangPmiMfjlhVaHhMu0VZbAT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XCLgkZAX+eoDv99KRMZHS8hRKd1tUXOHTP/KGoQlEw5+2IVi3AWTDCpKv+6X
m3+cU/UHNwDeBcItPOE3QWvd7CZ+wPS7NEYCssHqGYWdgwYd6jwp2j7bNA1o
1q2TIYi7+RX4T9WAL7a74nOG9KDxmP+k3R8PgKhO/v6KCG20ezY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZFrVmRiSk7O8QFg6bwRFIwC8PoeoJ20uNikV1KH2IuhfmFdJoJA6KYYOTadb
uEFDb1qmZVFjsJAKyrRVuTJpWoWawayo64TGSdhQiQ2wKvk1FaWNJr30ZlCO
UplFZc1r+tRc5AAlN8GPYZPr2ilLNPxpidKG/WAYicrM89ZqeTs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 90320)
`pragma protect data_block
gGCChGoN8iXfmN45E67wzjdVjDu/onCNQNyj9qAHYdgeEmBHg+Aam1jD9Unw
yEIQHZ/39amAy+J129lVHPp5J17HJdnUJ4by4enBdpLLQ8hAd8KKQgE+0Oyo
y1QbrnzIc7u1PGftdrmPeHfd3qh9TiXcH14+6hfmPVfvmhOumevy9+frFNHQ
xGDQSysm2blACrI5Q47A1kg6kGi7rXvJ8WYx2qKBsxFg/OOk8cxAnNxULjcq
uqbg0P0UtmpnnzzBZ24TzPUfREnjtGsxFbMxLCQjM4R0GTbWBusJb//w/qcy
hH8nMCZ7JXRVTa/MgGqHuvuiYNlTG5oE736SVHi/s4pX77LDATRhJ2fLyMAq
tMB2QCg+DeTvg0z76K0uM0zBJ+KONpa+AtCKILgG5N3R5IzVReQzVuKdYYap
n61zSnFBtwk+lPvEC/6p1R54lwstVEvN7LE01kKkMxfXEXZSSDzbskU4iEU9
xEaRaonZG2KMp34Ux5QtCpFhSgSY6LSd56Gx3eSSo1+YMlwW4da1aNyyiJp+
y7j3xYnkqgNx02wrxFekMSbD9BxPilAMala/GB8nqtPdcB8IfRgiqKRPaVa7
AK17wRqEyTRsPkc1p1cMWnAOuGxp2vERQjeI+DzPF/52b7ypCd0h5ANd0hTT
iZgteJp2I4hD4yBPT+S6I8D+NtL2vlLHaj5Cy6jmlIVWLp3lj8yHgdXyE32k
I3B6jOsl1TdClGrlY3uLigiZDNE4YwtLNL+LCjKHuO5tMSGFICZLqocKLiRt
l5ifFLW6+604u9NCcSVtnHMiApuQ9FFAM6XYeitUoKzZ+MRtOnEjODVYsPPo
VDx8+VEGaOUi+5E9+8upn8kzpkUoIMWZic0tFHBDTfwMxBnBYzAsaqhB/HMW
8GxUctV5Q5skBkKCAttPE44YXJ3NyvS0tYQ4HxBFJRSoGkpI+Gz/URAugMfA
3SLISaOiqZc4X3zLM0zLwePkD0CL9/B3Dya58frao+5gu8CdR2wdjp/cswAT
R7UVerrtrZTIaHdL3CXxypTCWMllmQ5yKw9AWku4Rc3XTF21vUVyY8UcLAM8
Q6LMLa0jD9hhngS69Jg/bywf/devK9D3rutyne1bfwBGWQrJMUfKDne3Mgfl
52MAm/2bpdRxSO+XLMTLQlGqvv5C579vE7fR98X4un2utGMne8rjZK/I+/jm
ODzJUVidxzbbAgB3GR9qJi7TpqrlYLgcBj2qegp4j3Bva1HrWFUhVOkvoz1s
x2dFbmJQ2g4Ta7E8+Q9q6V8uGd7owZvED9OsjqN3DKjLnmCcGgJW64/T6w9w
Pi07vJKKZsPIYjLa9Oz2tWJNF7zhrx+l96KBuIXob4Gx7Rh1yw5o4mxxquCd
exAw4u6AD9eJdjRxEDkuDZZw7HciXE0lwpc2YNs94C0Ek43UH8gv2KHaRVQ3
IhAuh1HPKJFFuuzxMU7ooDY1ScG/NEmb/m5qwxZSXAUvmj3+k3PrYOyoJkdC
Okds8viSW/eVsbeECtWE6ALCOslr0KbRb+qcRyEC+E7wBmNC09Sk9kTCJTrP
6+guvckG187eFx/fM/rNb7a+1NPTgPhN5NiMMjEK4NTCKiXio2RJhHosTYfe
XBUylYSte4iOkW94dFhJtC6fJZwvHMcLQ+DZCpzpE1bgeFrrND13YiPGYQPw
mHYzwEar1lObDeZm5OM/3HOMaHssrIjga3e/2O1xMLnfViRN1aejby64CFBu
63i87+SfAocAqMHnqyjAe4p1tuwF1jLmKGi+qomyepjYkbD5Pmh6FPXrpo8i
oTEb8cGngXG0V3n7AvtpoubMqRwPfOk2A/MLXcjkS85nYwZN8nzl2gvvD6ME
NBtWmQlYRMzCG2RuvUaoXsi1Ejjd3YCvjV1iVUDrXHHtCWsoPICziduA10Ab
tszmnVuEngudmNtGjS3prraGJdNIsj2xeHVG2jjKogqfH65VXlTBCycvjBDd
XqYT41e087PeS2MYldzjwrhfsIk+WR4Qad/xw/3IL5AzMAWt5dgaVHQeDYpu
cDllwwIOJtpt9xmgY6XA0JYbMg3qdPIJapmNNZpBmK9ddIwU4a+MrNuENiiT
hDYW/UYpwmyzLORp94hhcMmx+b2OS2AHJKy16aS/rqRhzxcZr8b86Zq3GRKj
wC4796wZt40PDPTW0YAtFR6GLVke166MHMOCRvRqn4mJYNqs7JyRzrrknibf
lOZ8L33Q9OmJlHOMy8w7dKvodFSbGzP4etOiXQ1NQc5p7iHPyipBm95lfJdm
I1b4fwC0wUXFhnseKRuWXV+jo2N1G/VrvQE6rsSZqXylLqNP+sqfIcvpsAn6
+SqDzLp1nk9jrkhwpzb2mX21krzc2OtLNA0P/gwEEwP9RMHdodo1s86jssnM
6K+Te/06XzCWvRhZeNSBEYEI12ut2CEx+IlzexCJTFy2tX7PeNwqxNFNYxmj
EQZE+N0OuVhah4Za9cofICc34JXsd8iW9hDpEHBTKonk9jT60Oj7VdvVSkyr
5IaPj1kFIuDq9chGWlm/slMS/9+oQovwBSp3Oq8MwmM4iPiQ3fXd5g9B9w7C
la12Ck9yEtKbJlOOp2gKxnzagjzCvxj+KPb30z0D8gEiXE+zWGqE+r9bbKws
wzhmPeIEqaNVCmz39CCQHkWcj96po0AtsNpFgq2FCZaJNvxPAz2+WLJ+m0P5
Fsg3z49IRWVkeYQkko62giggaCbJYf70HBTN5B7xOzjSLjMi2qFMnxTeHd8Y
LIaLqfO0DI1/9KlEg1OL9fp/JQjWCWf88OPwVRUrL33qdZMaXAk4Orfv2zSs
oldZoE/O/7fiekGjt9MlnHE7NEWew05OcEXUUBtHuNxlAh4D2W9b+Xj0zwHD
2YZmfT9w4NlDK8KqqvoMjFW0vTkZG51YXoP+tKGMz/28RPqPwNd5ADKJ0B7J
JzsSsBEfimotuUiROrBcFEZ68t8DumW/tLRZg0AortEpnD1r4XDKVnuKq0ze
G2T3Z6t8xCT4dvLQK02Jgs8lmgqAa5F8pbNQYMOyHfl6Qdj/kqjo60kLniZv
UZ5Q4XFQrpSAMGDHWIiO0f+jbSVOn98QPFQ8o4t76dp/PVKKRcCvoSxx+hqN
B7iDJxgko2M519w9FrarBbw18l+YrUxzvI6Z0ldaraM5nZ4MTFg4wBvV0UmZ
LQmn52XFt9rYlqe03A1EWs5mkTZjtPSUHxqJs9UaiYEDAlfPMDs2w/EVnbG8
UoqpL08IRy/ysyuiXL9Nma7P2OetnnbRp+9ANUb9R4tLv6OLnNRZZiJpGJ75
s61KV9O5pJPXLu3S/SJ8kowFAlpswShZem20R4z7rR3hApq3AbOKeZP6upPU
CXHU4SSgyeHKg1NrZVmqu3tMBeESkV8WyptVHKJV24vjoB+PNYGAzzagoXtm
CFAnxPg6L//ZwfPN67/Esg3qMCdUzMaNCYeMRQkCx74Y8V0jodQM/Kjrutis
wMXz/OSwtOygSRsMY/BJ8lGTN/JIgScKVDmtL7ftrKwcUCQsLEbh8li/Kpht
wQbuOX+N8KJHGOcFy4i2NqaTtdhwjHjkGhP4sr6lNE9t/ib3kiR61kGrXbU1
O/1vUv7UpkbUSKLzB8AdxnB4aOjyL+B849tCw3wIxPy2CFJRoGt4EiNJhr+K
x+os9WjioyvYUI/+at8SZY/ZZO/zq8W5UCHR8nXx+2S7ovl+EQnWIEwK53/7
TloacptgVqVEEWoEq0toYwt/AcjMqHA5pUQnkgoJJB9ETPyju1YHlijO9AAT
+4Ts+hA8O6ohz7+Osrfnqo98XIbz6MpBouKgyS0MN9fMfnIxuAe74OWYxWou
idST/O6dhtJgweZrsw5NY88TAmgjOORJag2AtAVTGkuxE4GMHN7LRnbF0OvF
pMQYSIFRV1Sz3ZfBJwH32VT9Dhsslz5/2C5wYLuJsLbsLTjahz/NwCCtAbiF
Yq2ZTTiu2s6ZPku9/2wRUJgkr2e6CQxzvsxI7tHfN0lJsKu0ydJeK8ifrpjX
gXIMvsbs4QVN9v1sZt0CTPc8kpzkGMA93awEKWwGjMkptYpSo1cmTTHtIrRL
oVDqTr8rW5b4yN06hVuoons4M6u0WlhM6+/a78a+EiAKcWD6SaOVnn86qLKT
1TF36sDMvRH3Z6rBSfoZ6+iGF745tenehFYr3ri3pVr4+BSdyzU0LVv/ChGL
7O1bQMVOMwsYqfYkJnF+1V+5fGuPybF3JbMO66GU7Bee0iVBl/e7tmpUz5f6
SyqEG7pSPD2iJdT/gGOcmmDMDIUFC0oeSG3masZuhVhTi3NA/0NB6awXxESM
YMU9Te0INEIeJcruxMw4xDm2lE8ssEbEw+hZLhGfs81zaggWsyUZkP0K0MSQ
sPqOtmZ/PCjf7GvFce1UgQB1DkGE6F26DdLUUUiAJh/+2CXBVN/qlZ3jzSq6
22xlqEWjfUF/ge7RVBAzjMEWQjJPE+LLcV9EHYeRl5E58hFD8bWXs2CXl+k+
1JVIH9kW2mKwn8yHTRXn5M87fFsguTvq18D6nbzJW5KLmxgNb1tjZlJHIFHq
DTsgYdVnWyui1AWtF1dA8UHIAWX86nUrUDYyoBMXCP5/p+X4PDHhTJKSCich
X1fSdz24MJwj63KWWOVtWztOkIr6z1T1zIOZznIFIu9YW6sOYgKR9JMNVWE1
N3Rix817rQDDgm1JrMsxik+xOvyCyxZLNpbPEe1Yl95cwLDymHm8HC63NgMq
EJst/5bXE7PGosRk7/QJoKr4DKRNA5y6ITZy+/nrNDiK4/CAGivzDqS3v28l
YtcK/xSH06aTf5ofdGQOMUM4MT0DfxtgPd7IOoSxeRLgHiXd9+WMmCsvwGH/
t9oq5kb+JOaaDMyXR+ivKHvpV1zFbsNyWdPdtqvSznO6oSGeLZ8FQMb7IabT
4bq0eack7oXqh4IOBLHwE5iC8TLqcC3bluTMl1LWPB6rnM3JdTrDFQCg9fMK
aTZvc9LhdrwXdHyY26x/iZ0luURTzdau9NFK2G5OYbLS4Z8IQ1gnZALSlt4s
DYPLweFfvD2gfqDR7HHe5K3X3Y845CopWECooOWyjHcjwnDQHMmLHdJjJPXc
J9pwV0alMtpN3JoaeIZj55GmXpDU7gLQuBrv7rsvGj+AY4UMFxVE24UVJVNz
K9nySXV/2DLxhhLuTXq71rX4FDFQnqpjdtkZGATOphjmwnnK5GPTVCYC/9hl
oKdPpXq+YTUO+4LKUL3tCv+QekbdXz0uUAf8qtvzl0M+xmeYhgx0LZAMm3Ai
zrAOgeVNxf6zklDjqjgQ7BrLWb1y2g/Wt3HuPxRCRXrj0xJ5Q4MKsHmfVYUy
TQ0uJFwjNCTzG2EAozZr2x/qc07NV5btpSw8t+2EGEgPfYHpP437CCV38WU9
U/9JwbIaR5BcSomJS+bL1idBfszbSf8gqaAn0k4Cx6nRHEh6paFD8YbllDWs
uxv75/MgsSIgFuPeCwa0saaCsP6l0B2jo4uY+8LF9fxnGJTPuh0L0AiIcLIs
nmYtKYYFt4ILsnjH417K5BZ9Q3rEyylUbtdx84IU+rsSfqHpDt2FM72eGW/v
Ala2jCqIabPMU6qwZmR985V/Pd8L1sOegwvRLNwJV48WX3MIAfXY2WbhHX0Z
eOJuf3j3q9iSyihkEwnimRCEejSwtlloRU77+cjER28HD+95KOazk/hJxgu3
aOj/PsNQ1JiWmq+IrZmuhWlcEiaBBnF5Ft/PFj7oUhniMknm/FkVEEgnZ8IS
N+M0E8JKLFBvH68pafUItntHQO4c8Wfs+D2H5IchdByzXdVDrinjBI3wXO4a
IA/6kDCAEhRJabgFiBblLAmwQdrn4gUja1YWQjfM3urmhgfsmXkqjTdcm94H
vGQ9FRMMOeV3lzKPNaGzLsVHIgOnPtZV3wSKnZjbJKDIRFRPza5+Y/CtHKj+
nTv9aUDDTPmJsYCXFTw1z/OnujETp1v1RERKOa6MEcxjwVD9YfpC7mK9eALT
4PexG1QBxEjAE9zBv/mgYQFpg2FmTJT1/Q8wW2xMdfHRP10PjWJ8Syetin2r
BwPgiBfE8zJMseEoArcfjRKZo5YMEj/cOLTLVmm29MENbQJhfpLYhVNel5xZ
BtOqXwgbfjr7t8zaSGolUHWOxw+S+pF1yjX9zC9T0UvQ21WKXUWi3lFD0VrM
HKWc6ZoV2qZbPZVldrsctNVMWSSxiSMNHs1bD8lqTbY1Qbdn7z68qwAjqoDK
JwHkyQbJgmBbzfGr2e8jKIrc7AVWeONUmJ6XMW+VUEL614TUsXHRjY605/TU
qVNCtWCp7u1vkgEVXccuIeZbFZl8nNvpcHdrOC/HXrjRmlF9HfD7OTt3/OeX
6stDsz907ct3MvqAq2Ky5AkGS39rdepq+5zfN3U8KmX23c4gCHSS94scSx9j
+QW+7qC8uT6cK8Po2KhEt8CsWFCqPI/GfCZOo2t5QU5XspsBI4rxE/gVqYvL
rogmyRfGQdDzz6ynRd6+3xa56cR6XMYbsGvE65Q1nAb0h0Toyb/wE/CaJIYj
w8V15Hq1f6HJsB9aT9bK6yaek/bYcNeUgpoJxkrbCVV4a0aB4rMs05ODsRcZ
YrThyQyyvkvB3687wE2VYQZp3TM2Btl1Jpvvf+4Q+dCO24JYltWVr+v482XP
QmVFqmwcE0bRiF3sYges6RoACHJHJYx8YD96eyKYOxpRiGehdBc1SMtEQol0
1AR9f6e6jLfWBSn5Zj28R7WjkBGXAQ9RJwr2xAcdmXwukdHxPoXuoiF0RdcF
iNSLtzSjNJyqNkvmRBgw9bXi3ERpYNcu1X3Kky4OY0tI+IOwTjcQ28naY7/A
eEwn9t8BtxlK4d2g0rE6+NhTJxwSennc6lZlkJT4HMryTaPuk17qTO2sUdkE
8/NtZ0oczuan/H177O7dMSX3L2T9wjZV9d2fzEDOG+1mCZRePBEprFP92Om7
FsrbOP3CyfnpKyvithkmWXCVQsGReK9ZPxW2Azgtea5Lr/jkts9kOlI6f45+
UFRcKERCJwuVi3DItei8n5SRX8/DhE9sQ8kB2UT6EQG4gnK8+SZp0+55qpaF
puAiRvggzONsnCSCECevUggx1JQyAgIeXwSHfLznEBViKul6P9TbjDhzd4cY
sGrRRP9XsNL64nXp0GTH0gYuvKKqh0ivQHqxeJZKVGo6BeK0M3ULICgccBqD
QjFKWO60L871x7NHprVBC+ybiwmSF4cmbAP0Ent1//tmKflCcO3pXtiqjI5F
I1CljdPtVROBfIFaefgM0XOZM8gUUvAR3fX+3bYtGG3Y9PQrwsXRyYKDWnP9
hgi2XbOK/sYUN0uQXYkaTzDkZ62RtH6Op4KtF8Mxd9IA9Qbwe6dqqZIuKVWK
Ye1t58tcQs3nVhwW8upmOJS8vX6Y15FgUGlR1e2NyqOS3vuiudycENgkClxB
0ugXbpOWQefjHfguintxGQupA/f7rbM1UG92pxk1W8Ce3gY5QBgpQVqMQAdd
gApnyHukc4S5UptJj3DudO97AYpF83IcIrrqSQsgDdCx+OWp5z89BLCaESQ1
8ej8BojC6ec9LREGnRtH+jeDyhZTzuoJkDoGKvVzMKDXQ2WuytyY+mT7/CYt
DbEEK3ZqqdRyZMZZ5LAuI5Wpl6k/LxcSYD+IaAQ8+RrT5dSjN3Hch3aZQVpv
BEA5G9xPfKNCAcfXTRZzeCk+f2dHA+ceCkkHp6Z/xDrRUEviScjTDc5RpTUs
v6UxfOIfxAQ6oLLkHqC3msHD9ZRRp7hZGywSjG7491ms+SR9DVZSE4l5UDxC
7Gz13paZi6kpTcOCpZAgSXigkhc6YfNsdQLEcI2nGRSr/m6zTRf3G7Duyv4L
aNyvo+xrv63FY5MuCSORXIaaEa05GEcKXAscSUghkOvZEePSX/cRQOx4t4qn
fRR15GC6ksf1sQmbL9O2ldPzne14Ig2jaLVicCWTRyB9t86Inq+m/FgfBD1Q
qCV01UuTvVdaguFl0a5pbSmJynlaIEi8aJ9emj5Qitp2H1Xtf7tUHomt8ARj
hK8igIEWhboOliM6ScrbBHtTHWZsxM08MBRge7aUhoySMav/VCpN0+LFb5to
eOUMO/uqnhjaL4OpRS5WgNJDNfRzpJbjCjcJTFs3cKXXTBpIovknrn5Hu9E4
1+p5+OJcyj52GGPSIRNubbfIDIdhZSLCkwN0p9kt5QjIiIpiArNxZurPxVOw
IsecMmza5vni2rHjhzJ48teRxufHkvEIYWSAvOP8mhO4mGDOyOhkVQLVgH8J
2J8sJjVNgluKbYWbexxQKl1TdSdEFfSuyj/MFmZFeSfaMqhLcTzkp1gUrJOM
oEgxYvAhDBtSEJ/6jERTmftCIlQYQ1UkcoPWhgcHh2LFU0fXjPTrm0imEAhB
X88D39+J0p22JmoD8uvH8TsTrFHCM3CugedZvsanlcYLN91Zp0MxIr5LgQK6
Vwj/HP8ItbmVoh7u7SpiDsr6y4dKdQNeMK6TFzR5103nB3JzdcHfFxa/BzM6
Xxcl5F8KNbWBeGi+shbQnOjauCqNGz429gcjEUHSyVo/er0ZHxgvYmNd9SdC
S2BK6+ers1YLTtLRHMFxvzXh00fzj3xa3PSxBNE3yEut1tuV5mDcvG+9kvT0
zBPamMV8Q1CVSMObnZbJz7XwQpj2Ge3ZygqIkkWN0SQlF+P27V2ez0Y94vkc
8vfWocWfaxzYEyqackxe0wl2tGdmxHzVn9tRIXUNAHCknvNt3sdOGTM18vz7
YHOmU4s1Dqe2Pz+XK6TvIdjjNTu7O7FV0jkLfZ3SoVUhhp4tM9NDEb+ueb9d
PiYwBtoahaIev3lrqh1AlxwCW1dSRGpKOWtH7HS0KP6WKf9QfuOxpj1KiZoC
3DgylnuZTZWMTdejb1f3QaUYfgWlXKOQQQvkiarFUeeP95/DcgsDn/vfchzz
zKjI3HOvjjMlZfnK7LhgTCFmF8iT98+/TFylzDA+inkdBI/oOoUr4hrDitY5
sgyM6W4z6eHaKrlZB4nrzKxviLuR257rIEkYdIjp8wrSnaTIOcU5Q7qPDpds
vo4aRbq+m08uOTY+16K8NXKTPONJ/QelCC4K9I6cbN6ZqVB3fyk8ujWTzTxS
8j/0LmI7NqfesezEpvh1kFU/EALX9Dz+kKixHLK5gP/FehGs0wVMATvMA+7F
TOjkOIx3Muu708mmVHKBx5afH9Nn5HfjJr+bM87RkOIntAYUhEDxxCB5Pm52
qJrACHBBJwDQAKxwRv307wdQ6ywv2O7rwHYTDeXqUsYdyt3mgej7FJXiSmz3
0itJn0JlUPzSRn3/JWPUv123Pl80Sr4DZ03IOzG7UafSEFF9ysr4YSsEwB5l
v+BJfqWZoG3nLgf3IwUOplaieSYKZTHz3jsfImfcIf4liot1edq0f9As09ow
UPvKjcbmW5hMzuY7o5sSntVPEjN6tGWUv7g1c0nt/YL5NmwxsRWo6pEwQf1e
UFJemiQBLjI7x/VD0ITepv/Rnn8N4qAUZ51/WAnhVmPzwwtJz7TQLlV6PNUt
wxx7PSM69++tPjmsyNFLVB0pxGVQSbJrA84ICVCjH2fwE6zgMLrqlmF7kzNI
KV5j/Y0m8MGJXKQeNCmulFOub6SH8xCtZxaVWK15gaZjU8JnSgDQurSWxZwo
AAQwFBU/uD7O4XuW2pp164ExvcI8ZJ3s+6e/U+mObhd+0y/LFkZPrYYHNLbU
zr5qntSBG035nfWshkM8KhvJmw88Ba8DPtSgCXSzARu9zBHhQL1sA8kc9LT1
ylVBoMgHnY9NNc63YgGkb5UoOkE+kxL0exN/gnm1RFKXqD4AcWcApt96ENMT
MUKcT21Ps79Y0s+i67APcOTqjkAvW4IRi1hj18bV3OmyIfqerbXIR3Jwy/nN
WOhK/JfYoP5LT4w412N4yGqNOyiOQz67MNaQElR3UH8AaLli/k/PaAz+oAbo
SGqYbiw1GMUUQ2VQKH4LZpX/Rum8ybaIVE18FyLLh2Dk3JQr/KTbCB9Ap8Ty
Yu0HMq5Grs9IFp0Vl9cTjOxE5UB+dshAl1Aiqqm/FPpD+aXuAhH91F8qymum
tqly1qTimgkwE/MQ/A4jLBwi1YaIrBJBvSbwBG7O5w/10QG4gmE5r1DkyR6v
ipx4SlHPhebOWK5OgOAYWb093nULj5AoQBMcv3mn2pkh8Exdy4eSi0GJYLyl
FM8tTG0t/LO+fbenp94aAMw4P/llSOECjZYExoC4HCgGvOeP025pJ//j7fOr
0SmHyRFhx1M7N/wmT4cuM5KXkytiO1AsxrSD52R7GPxBgCu8ysbRdxeU9UBo
AafX3vkQMgcvHAfLrCTxvtJN5C0XsqIats8PXLvSEVf+USgwrQCEGUpYHM0A
2b96EQunzRY/15u7ZMeRil8vQQolYhDP4I7YQCeQSoeNKUGvRCSXc5/gSrRW
03iYTFbIxmhVU+70iTuyMxjM8JtemJrq5i3unrQQNJs2YRxWZTX2PyCv0L/J
7EyWy62fbb/EePMlW27M9+ZYDVfeSwahy/1hj0VDCBR20KfJy7ZVKVwH8oBb
SBrxugKsBbQzuPJs0zgmY6mlkHYQxkGCW0+O6OUZlcwpVJ0Tj2VzbKqZBQCw
bD6OF5gPTsvj8Wc0KPvjPdIOUT4gKzU1lKMlbJCZdBNCyItDhYKrtAwY7l2P
N+lUgRLCpy7PsfYuSDgZFKti9MnS4+MSrDvPSniOOXcKgpAA/ysJXSs3IHt+
MuoFCRTvENysT09ggSClp+XFR0NZ0ByGjzDoY3Jlh290jrdWBJYvLVjHY/4f
c4lQdSAVXRbFIPz62WGZQmnbWRWOdXtYvT7AdbUlHQAdBANrZtXcQSox9MDX
DtYJbcIAMVduzCqRH6Zv9qiF5IlpxYPfayQlMODSPxovWb0vuiK/QDM3RLxZ
4g5UlRrY4QP16wV/smHFj7+4iAsI3Ky4pPfRi1iq7sa5FsFnG5UuaZXjTXMI
Dl9CfBW/SXe/ZZlcYlzdZbT/j658HGz55w2I1SDFfRpxaMa7NA54QBghwA6A
Gw+sQ+bfiAGkkeNkNPmEedh7q0NoDGIFILZkZFfJA4iZapJ9Okt3PCrOonQh
q1FIcDUXVhTftzKkWedate2AEmF0no43KGFq3Y31Hyg8T/joqwZH0JhoX1RG
XtzGjVc+jkZGte6ZNvRiiKvhPqunA/niDXBPwpJK5nMwP3E94bTRqHtQRAa0
BMViLsjL95D2Cu7Ll/WYxGdLfNCmCFk8RwQFJsg5+SiPYk7aEF322ctFizWv
ehEE3ACpIrIQY77vlSTsJHLbxU6XHN1GfjLB4s/HH9pe/V7Qq7GYzPeaKSLm
+uSXwgP6QW2T8E7mtsb5Svc07mRGMhjj7kyMGJ6qFdM8Wu1cnKyaTVKXF05d
7UDFbpG1stRNEhE3mIh+fCdExkgSxvZM7fRfhoceOxL/IRYcEToKpo/DjL2T
L6yMSU0B5NcuDhHRB+x1eN5Q4Lop4K1cYQtkA7BAywAlZFpL+y1r8X37kytO
Hy5RWV8Vn05zEgFONUcYaqNn/A/VfcefFFXMz+7Y7Y6BspyVwPaViDqqX6ce
VrCdKmwBa2AkbgN+bwR+BdMMSjHWo9H+crV+n9EstdBxhxqYKYfkuzJHiUx5
he/hde42jtUmCbvtKP5oUa3JJjxSdXg9HqamrlSRjkIEUmc2iRTUF2CT8KP/
hhaaLe1WkzCv9cEsZMVn0pfLajl/sFxVYV7qqed52TRUJyyqoNwCzYb7M9yD
7/nKmA844do6mMy2LWu8UpqzitMY/6u/vYDKqxgNBoMV18X4piz7J1IW+YfK
wP80f1PGoRJIfUvyYaBiqh12TSwctxT2eBOrk2oBoAdreOv5ihtpt7W2s6t6
fyJkDsdtNTJvzIAd+qc8QGpTTycIveEfuK0h2XYx/VX2+H5Nt7w8bcleB9HO
ZZhEUEEwtmh/BkMuoSBObZamT8wX6P+eaJTkm5mXQeRqekV84PqNGQKSJ8LC
VaSba4Tj4jDD9HlULdYiu2wX9JUwKDgd7D3tOhA2vwTJnL34ArI71P+KapTA
Dra8wbyZ/GOSW7BSkvf7nbJEWKq/jFmDl3D/sPi00380rM/YchAVLA83El/6
LgrrgXy7Fic1Z9aGEfkfM/C92iSanKyfu//Ym9fy0U5ltIB/5t4VMKeQyBS8
/Z3dr7sPZOJC1Ouxg+rb7/ShMJweWHUFx7S40AeWnKGjxTREhiIDRMIVwYLy
+cjGhzRfNk3EOyGkJmMwbA/JH3TeaX1JW4r18n9n+xpknKmlkl0gMDzQ/mru
uZ9B0dhmMwLzrH7yyB5mEFJZfs3RKrM/8TFcsy93uCryFZdvQB3bfUlBGnnh
yWp/F+BX4EZAUPdalMB/4wYkVw9ueNcitMzYctNWwK8vMmoR1+sFg6P3VnLr
gNSf99FOAI1PZACtZ9+oKSUJyXDUTKpKpXdv+0N2evpWb0+z9H1Z193hOFvq
Mc2pAMR6DbyRctPjRN2slhUaCHJyp+nFzf9m9bpcDzLcw5yxCSYts9Kr1tLb
TyGi2ilunZ5Z92Cir0HdycPVNzF3GuyHTcqocQmSJp6SvpcTir0T6XtGEilQ
oRtfy9d84ZbiKtRvpmmbtyxzS/m62d5fOguzMMAQtPQB0pQcG32XFlX3r8+T
RMKt28nHRJ6Cwyk7C7WIMzkp5UP41sWLolfCagQTXF8BnLq9+8FOqQqp9lyr
Ic8d4Fr5eZZq3PjALVtRaxhxDYvj5Oa9EJNiTA+fXYIbyJ9zLXEHRI0zx1Cr
r8njStG5jiU5fPn7IunXRBv6lrLpmJMjqjeJwJbvKVdS6NDPHMcCCrCqfv8j
R+PjL3VnmQ7ULZfdfl/hDcVRKZd1+kuLTKEaK1lahOGCHz5qiexdYLzDU6w5
ekP2ZT0lAYC5TlWithpqZYSzMnmGeCYOwr0chpVU+1CID7qYzNNUgzEDs15k
5y/bEZhGLc2idOUoefkZO8LbTnND2W9JyNOnH9xagHpquX2vWdpa4vbHro2x
/ft8AockW/0I21vQxVFKMOqZODHkADreMQOSwNI1M0IqADsN3Ot0yQEypvOr
mR36pVrSpQHVO5Meb4j0M6K5n1s46KmLOXykuG4tGlKFxz6ExgOwQRA+VWdH
pwhy4o6hHSL4xTC5lKzbWVcPnrAVpvZrkhA3p8rP5RLDQlAQvhsPbGb2pLCo
3AbzqEtLRSX78DqJnoGRqMbzvEjW0S/rfhUJeYRmZkFBM8P1aeECtUyP1SWz
M5p6cBDA/B46FPg8vkTTF04n5VJMyL6QL2tN2zSKJP6dMVUcj+M4b1PFbMF8
r7ccY4zyds2NXa3TsNHQ+JR7+UJBtJO6XEc3l+taZtnYoYdZempFPJBHk9pw
uR/wqO7COSX6tLa/Qk9V51whxUREWlqdaqo8uEp5Yaxy8OR04QWY4quciMhF
YhGHzRNMz5xLlzXc8o1Ef1BrU8vFG5FsCDgN9WebG2ayNIgL37XeSyngE7P5
EPJmG3aqJgT4g1GOXnTea+iqx20XQC9K+o8heKh8HHZyiEire1uJ2d3MM1Sn
k/NJh0fuQzIcJt3BXCShWimEnrZrX2od241xNBh0Ced2g5MkqF1swfa7wZW2
lI1CDKxlDL4Wn6DOlDZyRv6itOdCcPSz9SyATggkKNqvMMVnoiTKRh/rJQHw
g7IHRHPO2eDKOGIP6ILPwvJWwSfnHwwOaV0YTG4sdzTLDXfu41jR7tmtepDa
cLYM3e8juZAkJdxD1h75Myzo6aYkKLd6p022cB82/l+W3CR89ZMZw3rI8NKk
MYWv14XFk3xWWVNk3fm1jypzgJMuCeA1vj/SiDSHEqNqatB/4C6GWEs+H2Bt
pFGcsA15QPTpTVX6H2bo6aYRgw/brZP0WgI3ZfksqSD36IoheyapuHTOsboK
wHlGppNrp7Etp9cPSV4pSJ3pHRkLbRUiZxeBpkA5G1bBYaAHwRXlBKaYumVK
Fm0rLAXVq+jKlBiCUgzbvpL5kzl8bxnth205WrM1XbWO8mAcCvJCWAS7y0RF
6MeHk3twymE5jNoRR4p16GGIii2NAyt7i11KE6lr0gam2FAmDNZe3cWMiKlf
i4M3HrTLC45gDZyR+5OiRjVnqOljOugjNZ3BWFNRif+H3GFabkIu+J/VEBgp
E1GJywydL1R8w5qRnARg0v15SRjiFlXYPTaa1cuEwg8CxeCBTiE0sMqwbe/3
so0C4y2WPDGhpWsLRlBPsSHK6v6jlopsh9zJoP8+jitcMWe+o35ZPJ2tmsfI
VhC4myKjVWdm93rDfo6FGvEUqtS0oW7qszYPcOvUETy0DPW0qCujg92fL+Rj
28OOMxP2ZqObi4TuLoJ1gDp6d1tIiJ+I6g9VjSDksionUJJtkljkkR6v7Im6
1wYzeboOOs5g3LXhmwmfMotryEuU1TTiEV3yrypf0ZxyH3MJ84LtR5WYDNBN
+wDAtBXCru6VWbm4MKUyK9JfXTnaHBTb7TrmamQStw431evxQa20Sk8TzRTt
mSOdK42i8TcBxTeOvrMuefFE40vJro5W7A09oHdOcqPKNNzDpwoHfJlBkQ/6
sGnHKkLKWg1VN7ks5r8EJ9D/70S/WygTBidK467MdDrDiKPqwFrUukfxoHxr
5AjkNra63eRZQZhMNnSp8Cjq1SnkqylKhWJ6Yb2jSx8OTSdEZY8zkQClRy1L
tJbLYECKyxIWRy01p4WYYVIIljcQMSX4jplGxOQ+HFxixaLb7FEKEl8wIhuN
kpFuWRs6JE2WaAlCbs2a5TIwHT4sV/HGBq9Q/lpLH16SPDg1q7tEprX9moln
YCi/UZ2Uqviesv3PgJoAmLbB+wWPIKNFGcpVLDqSJCqo4Rn7YP8FG8c0Mhf3
/vULWSG737F1B6CBkxlJYf6l1ioILqjZqMEJyLoXejOXQTrzRuwVGZ8t0ltv
rkr7G/bfeYVcfvudW0KHygLG623LqFtUaB9lPlUbTgXr+2wxVeRhaWtsNlDq
Kb3KDJoYQQy7ElnBejGDLjgC8cHmls9xSau8L2VxFm89eiBO0R7TVqACWu6D
4fJAKStKBAlRnV46stUFqaRMgaodxmCDuqcatKjvAwL2ue/vWyz/XwKamfnU
EpXXx4y6D+OS+KSALwtlLhwSlu1mvaiHoPqJpY0mw7Xf92AdwCa8ZORrhJmn
mAAC7E2J1H/ZCvOB4g8MelrBoYd6lYiY4te1myioyAsRDNkdIGwPjBQriK1u
kvy/EQHIqWFvLsKWyBgqx/Jb9a34H+djb0m+DjcVlkGgbkuO0R2ckLNvakyW
TBcWxJMeDdQkoOMtMOBbvkoj+RuRb5AucsEnckD7en9+tktvmfRgWYM2k/CU
W2ixW8Q1QwfPYaEjyOYs0kTPG9sTzDBkwS4IQmXFW+o1We26maWgLj+qZorm
hgwS6nkgNl3wvpB/RNijfj+utNdztdQL70PEDo5z3qAeevC/Ta4zKnzha63H
d056Qd0GLGN1SjBjd30Ov//Q3uD3504rdZAhOI/XXXDbqjGIIzKOn2n9ZEWC
MhyEopM5mskSl6S9TRgjcaGqg4MWLxurUhMFAtrhoavYU4GzprZPfhM/Wcrt
31c52/VwTwafWd4/mjjT/X3PrVEmo1cWqh8V3W7AW8nMi4bqBsTDek8UqOVB
IFq6JP57ssT/HIe95KJ3b1DoLe0KQyDTG8IcUtmmMjnXSnYspzu9tlgu6tC8
mWK5T+bKDC6edZHjEPe6wzHCQLnAYG+pEvCnv1hc8OHgV6UEA+Cl/ysFXJ5b
Nn+mFCZidux69GeoufdGiC8+57Cl8+mY6YZPZb4xAkf0zMbMTV+69LaRXuYS
5eVKS1Fmrjf8OG25svDOOBowIXW9d+6fckD94L/PbsAgTnPZI4aNIQt4zfNi
7DxDvVM6RFSqNNBIFg3r1cCnJsTj9mNI7RGqKi8ROXO8VSGcv8ZhDEIRcQFO
4ORAMfiqlPKndACfXTpVgAoBbKp4ODqUJ4BQh1NbBXoxTXIepkrwNpOMByph
bDlFYaOBkgEKaMuJ3jWPttVSbV5dLa4O4vxrI6R8NvIdLQpOIedwG+1ky1RG
hcNGvK8HJOxot/JFacgrDAlYHVSINeqRakV0kub6CVA0WGlXEM2T30Up+aMY
D9f1VGZvnHHsC0bOyLhh72nsrGsA1f5hHv8q8mhY0erUz7v1zVDNbYJB3V5U
6ooFGxKEFFhgKXx62rL4F2A8xPseU/jpnpyk5b27OzHHLgR5n0Qc+P0822ts
9w72qzOThYpyGYraTzH3w+UMSYDlEwinCKLOloB79MToPwqyaCJGuo+ABlct
EzoLgSTqVm1tayB98vmb/0usQefIwlqz0+LSX/31ibnlG9zrRGUNd6+ljOET
c2nATg+KZTIH7e2k3/cQba/Oqvc81vW1diEP79wsr4KGlHJOcmqMETDut5iI
kf+iozle8vYyzhiqOXkwBBdi6gDJ9fWRkrG3ICFy0oyjmHzG62e6xnaakrgL
F40uLulqm0eh1OM8LUvLiqiJrKWp3C3dlxeZUKAqtFtC8qTl1yJ2kbJ8M2RQ
I/1cLzO639YjqkMHhs3y61wy384DAzr1AXJ5lXNWl5PI7OJ0O/DC/95curPI
pa3WkSEa2qhcFd5YOhDYdrxI+fcV4TxmaG6ojb634CeJYfGlbZog42I2UGrf
isdm0iqsx83F7RdFhd5ugd2gptE6I/DV/pLuQICPb7dqlM58Lt52g9DZSevX
j/irVHKVQebW8Uoi9zHbsZDJ4pg6Ns1Ak3/UvLnpdW+xD/fuDMw5usagxum/
c7cZnFAn2JhAF9luLGo+TYLzVy3cN2GkI/bcrOHk7Fpx9oC0jB1cxoxRqpG2
u0tX0sPdcUDGfFDtyDzM62qKe1FEahkFzjplBiEnFehRHrvq12V1ALStNr9s
lQOiEiTabQYyb9tvMohhvF9Uv0Aaoqf/HuAjgfNnHNI34RvFuNWy9581YMcd
e1yp6R7ZR9/9jMv0QIXmZT46wNhC0Krl2rNZVip8MjQ5Su9nROmL3Wqha/+/
z1Ap/YNX/+6jCT3n4SRbUEQLKliOa6VTlrr/39QsDC2+Va1anp8bMNp7hwNA
g7ruCAlcE097WoXdbyHdUsJx0xOZaYgPbvbbifhlgGDpLFII4tLaT0A/iFaJ
G4X5U0ffibAH33kJ9K9G7sRTXpqA8JpSUlxqBh/qikpVyVe5vFHzsq5T8tN+
SGat7sE0gY4K7MAGGwBoRcGj/5f2KD2+zA1X0kIyxGB3GlzYgZwb31kiNIFw
0MiMg7OQhKcp5vBzJqB2/rJ8qeSTb2dB2AdWajngnRr9a6cxyKQcdra7VbtR
EZxqj4+xzWBvsWJ9C3/MkRpBOZtkkH554qv3ctQ1aAOZwT1cLLMVWYkZVnen
r9boMBSuCkNZB6GRljSy1SZ50dqV3B9pAGwxlZlAYKfKo4Q5GGvYYXcfxqXa
rynwWK0+SLwShk2wbC/KMhmjg/Lebe8KdnWJpGNhMXMKOK3yYAtR1Hz5R/F3
2u5xlPEKj1gWW20yyEBZBi4MaIsupjCgD9tIzR3MNInBI7EvnbVHRD7LNdMP
b1z//CJT3OOwVat2s9/PkaF2cCFx9d1PttpQaKwwLRJMmKconc+YfwxZXen+
3P8lHa1sTV9Nh4mVviEyQSX72z4tIhlkXzDEXVuTjaPLpEPoHGfvLUZQXfFE
V6bbcNrEghXrnpyfGvhcKyU5pmcPzGUZablxwE94mod43bx080KgCyXm5p8u
kLMXiK/UXQgijwDFFr9Vj5YCCgPhvQws5ui8jwqUKB2pFvEug0zBXuQZr+2W
jfJ9Rj8PEozgfjFeNB6evUslFeKIJugJo0Cxo/7ArLcOaryVTSbqVuxd/n/x
5RXlMSE+76oRSpYkRD/VN8uPyUtydrE8wCK9+nLh5/A411rD+oYxPQIRArcG
u00lXgKMoi5LWlUKRBIzB8uI/r03QPx2TPZzs5l+EO3iY0TgLEHTSPoE5JhC
qEVYljEdeJxmoCWyrnLcmrgK05c+VvRDGX0Yur7rpnKtMA75G0riy6LuhtUL
GYXUk1b3zFwZsgqfzGT3bTSV7h7ASZcHpDz3QLs44IDjFno6kDr+7+u2RbY9
e7KlPH+1RcBmauur79DsLSYvmQKAXfur8pL6Pk3NJUxtpAhjjbGtGv8lhX1I
52FjZatKr1Y4YNYusgYTyLKNyxjP2wfc4WM8a0xtSG4Yv4IyKjlfOzvbB9h5
lQoWHTiqlckCrcXMyepkNKXsnVx9fuzyxV+B+HXzlDhZ/tAaL7uYchXDqvEO
KhYVZeKJx29POqkQUh7Iru6t7IKg8i8Euu6fNfwa83rQ6tcqNNzip0A+CmfZ
tkENbxe0hW0HTr16rkxg+NMr0zDhMQ9W0MBsAko1ydzHV7e1mCD+p79jFW4O
qZmROkiGbFDcc0wtMk4liLEBbpOfpnNxyO5NnPo3rleC/yaIGoCYfZO0tS+Q
DdQ3rGE7q8PIrJumb/pa/AWOwag1vCEo6W9if9BbOEhSvyWj9NoLHN+U7mWv
Eq9PgZttNWg+/4NX2h1wdkmZLO3zdejuqgOUl5JZ7ql5R7gx52uoXl6tmJCw
sSBITauEgz1DS4qvNW2++RCG860yjy+iX8dWHW3iCZgFxiKHsqbfh1YBjWb/
4OCiRHPTlZeVNktAJ4B4F4BrRVYTB1/HwISp8wxpd7Hy0vTkbv7imI4Y6DuC
k3fGhDABDp+iioFOdbvIaTLXbWl6SZ/3AT1a9fflyCV7O1bLgLlJd50yFN+Y
2hvPLxVZAJN9CPwU/RcrgdddC0bSV6ZZXwUN5Jyp3Y0mTCoaMxtrIhSPzpoM
R48OF+SLRduqucceJUYcQ5iZJsOVqr4yLvdjgWruBHisTXRzxT+PLipUHIAK
/SrIabdbKY/aj65iqWgkUVZVPHEvqe/qFK3o3k0qxM2hVDEcLMDaaCbgb9ae
fVFbZNaAnHZwbHMq19ctB8iYfUSmcx2QgHEso8aH9xqQiRCiYRv4+8ZuKrJs
wEGQx8pfYs5K4jF3wu/cfWA9dFZYGVCfsvLVABKmjW0BgeamRvglagTfQOW6
LkioYuz9acqGq20mEC++XyeQBn17W6G5YSROFVJ0zdkVY0PtnBM+vm45PWSy
gQcYxRNxroO1Gp4lw60+f/hqRXcQf9kcX5pJSR2uEiuQcmC2N6awYAPPodjP
Lb/2ziqBvxpHa8hNnwVJUpknx2ny/pNm2P3qRys8jhLSzkwqShc5ie4n7+5n
TaDniLitZqOzWqRwYyu9rxKW/9aarh5Yk/xL10kCo0ATv2QOXHtHgi8Lx05q
BLvunW3j8B2PsvDqXwWv5aQHlsRv5RPUJYgQosxXwVd+1ANQXLOHjQIqX0gG
OsEbs5WTHGe3SdtaJFOG+fT5Zn/3qFRe/v7uZ438iOhWidUZli8f+MWeFTJH
PcVlZqvCXLmyhm246FuZNWRpITrIoPdHBMXFyekGk1tyHVFqDFagE4HYPjWw
lVuzFY4ro2YkLXAxJ3aAhmwqw39AFgGqgAtP2fY4egQKT1Dhc1qZmT9517z6
0/JwWADEIDUQ/G8qfZGHQuo10SbJQPnsfiKhvxspZSlyj8vdQp29Lp5+7KnX
1ZVrXSs6ci849TkKHzUKKHG1LZmti6X1bNNpYCWFwfeV8ddKJc1stAsooef5
uNetpbftYCVh8Cv07MDjlYn3AHQVvw5R/vlinUX2F2wSyXZRBd5V89X+W8yM
j3RsdTnbgcP7/ukQGAeIZ209zIMJPoil64kNjHsDn7BnzCdcNqN1+Yc3+qs6
slIHysa02MoMikqXxIRHg6DfNgnoaUkc78VVB+03URMsl5o3po4p1zPuN4p2
ow04zHwJiscl2g1dclxaxxmJyA3Tcw+i8J3lsKi9LaVPXHrCHyIKqXxYW8eV
aSBQXdMKQQqI9Tusf+w27+VhhRl8WRF7GZV9VjWODCcw2lNd7xcK8zcCwmWL
nYMLwsAuX2+zESo+sDkTTrzQqogx1TbHY7hS2XyywkdW9ZVGqfjfAo0811zB
TyWFeNjg7GG75DEXWPYk+RrboycevYwniUb+IfS7Maqf4WCzMiFM8FMrSJEe
LG2Y6tSxUwCMVnilnIkMYxZh1Kp+bRNuMw6VUOOkv9fKVNFhvXoiNLqkaj3N
m8qvCLZKipgz+g/vf6a6jw4s3XqEwUWUdWlHvQFsTOBfZwZafyn/7WGQRKG7
czDvv1sYmXtIsJrsa8eik1mKlOZzoQGTYqDudHXAibSob29WTDeZaMKlq5tt
44zs9LwvW6LFMsLx6IoltnVy2TaGZ+CR2ifeaLQtf9K0bHMcnf9sZmksg/2S
e4PcQKKuLHSUguKqVc7mjN2z79z9kqRd2E2ONk/fP3s37YCDzWkmbcCxnS4F
GHM354FILCWgQKqyLxeVmK6kT5mYR6PO0QPNmC3trtN11PjEEvKXLwfiYlUC
uTIZ6FWrCTm/rB3/qHAoC5gNugtjgKjFvJ8MetFPm5pzT5IuiIFPLk7XAWAx
r+HGp8XSf7N5vUI6OJFwtijA6KnQFhde0KpD8cLmKROeGwsJG+hDRpUbhsKQ
IzEmFtt0jGbYQZzKAXwhbIAsfQ9FBMsTVKo5DLUT3GfahAemRyc9A/H4dFlU
PSSVchLgs0S0f0k6igGm7VJes880Lh54Auook43BUeica37XQbyiVDql7g9q
PyNUWKLa/FB1sROzBdnNu1ipEkTbJshRZ8TlYkU4llron9m+fQoSHHGSvvZK
0vC4FI/YelKuaQgGzGsscR0EfKfSgiRwhjEFX2tncjKbuOZIHSDX6WbN0bCE
7Bh+o7NtnuAnNc7KwjGls8hbQJDH1z0e2aiQsAQQNjvOcDib6K1JxbIjasG3
f9kNHX+2m/tMgGgPbYbjG8jld5ofWjCzBTunz5znxJ/o5x4WLfHHvhR2gY92
o/rlfxcsdTrv8WV6/fVhVTSPCsXSS60pmorlNJCnMxgyX0+pVpsF1fTRzXo6
XesYIjrRuj6QuisaKxWpmZYBkjDyuGIFBQgFT3bVH5rB/ZuuIpNRzWixzgRy
hcnFAIxdr5Bhh2nF49P7vHFsscsOtMdTIJghFqI3sKQtY0KbzbiTGGT8n+n8
Qbxkhtqt3HGOH/8NtWZ+IxQMYlcx0Zjmgxhxt1AN9hGT/zOVpluAMWveR1zc
U5BCTgzEg14Fpy3QSpo20ZxVCAzPs4EUDkHqkdpuFd9xb5MlAniYW2umfGlE
/sE3ABeTRg8P8UPg7f5hn98twqEMxd0TxGqggtWXDR1SOHl1ujc/fcfXxZd6
/QM1QrBbH4DfDAT8iU70mRP+DW89mrxhrV53EqNvqfFARZydoQYAjkyYPSr1
BYQ1p2nU6Wjt84+t+5TiCpNHl/w3PVBrRxyYKt6yS3MbcPk9pGw9Xl6Qh+EK
pK+/lK4JlPcyLrxzKs11TebWwjlcLV6XoDJ13SpS5pEr2t5IROK+FGMzWNok
VtX9ZQxivG4RTGcy3mWTNh7B42Ay2WlcoEG9qBxtz0FsVM+NLjuJDECJi8tK
nWfhEsMZ2wsvty5PQvojF7hOG06DfXaCt0QnG4C0qOYnxzZ67IzpIHiS8CB/
9mU9SiSnNcFhe7VXbnR0wUX53PgABGx/iYtbZDv96SxAR8g3jQC+Cdy0Ha35
ZCRwE0TK8hdoFeLWX17dUX0h+h52PHKDttrV72cj43G2EusPTGj9iWTgxD7B
vn6exmtVAYbq0s/DdHAIAsaXMYkBJl0ZKNk6Wu2Fj6L/OKfHYHmrui+FFUpK
VK39biav7Tq7V51Al9TlYITLlkwWCSy+ElqOGxUrgr4pHUJ76y3umAEA+pov
y/e3RA9u0OgDfe6yroaaDlQoeNodHCXH8eYsmZ/vubvsHSxbI5BgJ51KaIeZ
p6o0HRhadbxLiy4zvf6PNDGATUh5BG2Cdelu056QJxb0tLslgKGOFyW7PSJn
CCvtgAaQ434pl/Wk8+CM+D8EoQdA+4ZKgZKWtQ9QOblnOjXrFoN5Xf50RKfX
T9wkEPxgI8GKoGB0SzOL+6Tnh6fqHOryQwTqVlpjgKZWQ3ezEaYU1FU4KK8g
VmhXu28eK2bBWq+UW9wSbgQZGvOW8746c0Ck52wwkvev+CDbBxLnieAuvA7Y
xbaCIBn8r48r+aYALvInQzst+0nHKSjWajpdteiIHWGNAZ85FxLfFbYy1e12
Wuii9nxT+q3v2dZhbZixPDS+Bn/nvS0iw3dODN19Grb1arCk0yTkV48ZTRT6
XH1AMQw4za7ylpbsV+1Ljxk/Hxse02cSyOUvLIiKVd0tJY1Pnck1BuENY10R
SPyBDSXljbwstJgCQRIO1c5OnFka4W/ix0MFMl1i+AjlYvnTI4uQSeXW4hEp
e+nFGFRUHd6++T0mt/5lbsO9jEphg9TabkOVzGhs0ZXkUpi4NcT3NsSpgWIz
C/7zx/l3JY9/3IIk/YrhRqSIznimChoadYkg7UyIxhjx2KRVZHs8v/IxYv/Y
Pum1MM9TTGAY+aWXTVWJY138qfXjDM1P92+3hGUBhf34zshlwUhV5M8jsU/A
PvFiFOmi8ch2s7oOUITxUPJznhr9DnoEr70cnVJqc8cLA0PSVMn8FjNMBEbY
0TzoHW9toc6SKX6k2wDH+C2+K8yOkIOPs6V0zP/H+jq6lI7XtfhKKvyYgXZA
FPOn8kfL1ViimbzBqoTxCR52a3rOIcMqWOUCRYtNCgjf4cpxc4OqmyNZgo5c
BmOj2wy//+dKPXJ0KoQ8erN+aoEZPxLhykPpkJF51TQ8o203RTWomPkmUIPw
B1fbDxHSiEUDg7Y7OrDJBnJbYUcTPc0ZCoSd2G+QMnp+CqVjArWDxO+RJpkA
flWP2njBjxZQy/Mc2efXYVqg8+eK82vLEW1aJX8onMvDMXVDYHmSWdXbm9xk
Mha/ILxd6i7F1vsEuTalq7xi1ORHCuqNwZKEIFt+7i88iGtGLmuaNbriaWJM
Xqj9xSRm+C4LhGs2DUoCdtFCxQJvyBLPNuRY/cQtMRmaZ5D1DjyR3WBxAyFI
xVtnj1mrJh86y4DW3k9c21wdlht16Fsb3Fr2NPZlpgA52dzsZQWkd32m0959
jDXlxKSRVbjjCbY7bkrM5Xgqrh6+qZ6d0Qf591Dkoihx1Pn7XZmsgm/diZz2
mgmX1H6LkBSnObKJSaUBriU9MqRaI8sALjJw45gKFfeOWXHHZI0HiyAICWbX
i4VNPgJXQxLaWCwhsoKP6cuW80kqOsM92+YWLzYxnDLmDTq30WoGBlwVKOov
sbpJkf/wGkIvQOhe9UPcRVzXqhvLADmdQnC8FRKTXtNf1KgYHx8QaCkqiMir
N8sTPaF6PWV6lG9Xq3ZxRybQ4T2GFz1uZG+Ra+f6nE31+NCwe/GphoUXfqPJ
Biix5mi5R7RZX2mmLPRnYG/aiP2hLaBZyopR7Ododnhr2QT40FTU7Z6Cm2s6
pr8NySpgi7BgcMRtacneBRZnsoLW56dVpPQwp4BDRZLdneaf7T5VxRbfnRwZ
R0O2su/WKxZJIFIdavA3v6O/g3NlpmttDsI/o/PCEmZZ9Wvy3Imjh+GpS88U
slG4aRGIVofadCQCVbijtMuTMErFIJhmv9YO5/Uhnpa44ZI298uKI5H4EdFl
lFg7a5Wd5PCXHI9tHQZ/Q1RwESZj1uL1Q93OQmu8/VOfVy5+HLYs9J4Lb7xr
Acga/QioqEquUucCQh8V7i5L6oz4Y/Ef/yvmmQfCT0exR0B/AA+L5+owCE3I
1vpJiNb2US+Mk7xB9+1ksQGOsVeIYfvW6G6Njkm1do/72W4qyyykmvC02be5
fYx5Ivmbg5+T/4WLqY8GWLMUeALPJznr0GbvvFI31CnM9TJPugEX1Z1oNVw2
RRdSn4FYhkjAb6cma+jxGREx75RmTBCay57mlLcfL2sNonfgXOA66ezCHIZG
LWe6qfDE04zmT9JnM+0yacICIm+6sqpnU+7DCkxZs1JYpzXLZg35akBJ1Uxt
kKPExv96ngD8tjPpfj3Xi2wUjnGV+RWb2bZdCfVg6jB8QA+DRYDHcrObDOwo
VspjHH73OciS503a9+sFf/IK8wt1whmmWiVAZUDr2pTRK95x33+6wlh4DtBs
HibwkdaDrnyU9/J95Wj3HMXNzMO5jGcabm1cpIfkH2c+FybF7+mjYSE2beY/
t4unPPckwPRUNxP12g3KLio6tMsAghky0VA/pHNaIN+GjN/xpfhVD3TLRyGS
dGpASZ0fyATy/Th0cJaObPWEbM3DSBYtF6SP/Ibqu1+zmFnpsYbjUiK0SyNT
xGuxsCCFJ8l/7g3FyVPUzMkogGWa/zjPa4jl2b7Z6ZjI701j9bOvBWH8EwYP
XaTcMIB23KzVPU/NkE51dLBUdQFFI/pIb/vmjqMoJsa48Wh72+Qr5Q7Pg6v/
7DiUkf15VXA4+6hfaUj5+3zwiupkOAGY685dpqzrKxQLvkoa4ZRt1PoH2JRq
fmr12pgt3TfHaNab3Xz2dxJli3SOlGqSxRkcc6+KpdRYZvxWGEGa0NjXdw2S
6X4PsJyMpnSsL/qJNWT0AFbfVOWa7fcMtgOY0/KESVO/RE25ZtQaX8VnYmjp
t1hMUeQvQ0YIXmQBttMzJcQ9t2Z2sBUkJ5NwURU3ozBwE527qeF3UV2UNUzo
Pq0m7gdrDpEN2Wrn1JUEsGxqeqJOI/WBOSRsnwZBvYToWc3o0DQHeflfz7K/
tGlC6jnOBzLn9HcEt7P7CexRD7gdrgIAFRjnCpVEht7BwiRrddNEi6U/VTz1
51hdUEau9ZFE8fLFr1DHjgsmdGgFs6xKdNjH3yRROTO5Hnk/9UMkpgaYpeIS
WKFdYNlxlJCLYAOCS+pNK7SOCmsFj8/jtEzvdT7i0qKDCFaQYi+jDOaQMTUR
NBgYxXo+SbXl+2wYKIj6WS01Bl/H1CBFkqBQeSJpOuGa0y/jT8RSarSWpCuJ
9RY0uP4D7NEZtxCu/LGFeAQOfbDS4d0b562GcZ2Alhi2ZLu2DYbqGdSf52bN
SCfH+lsBh+uwoHetkVqg99XplxCfIycaHvoHc2pRx0nJIoU4eLHzr4p1SFmP
/sAp8Es+lX1bn7HOaPmeVuySfusglbNcZE+0qaMtyjaM7Ol/+Jj+NL5eqc5D
rR/CEOtUZF9wWfJpLz+3HBGV1LE/KEPBeXCTEFrjNvbDawl5r+mcbLP47WqX
Lx0RoFLS+fr3zlntHoVmpQRxt062LX8DjdzRL5rRJ9j+J+IveEYI+neBxGNu
B8CE520LCekct5Ye5p/F8qKLsiO98dbmruJRXjjI32NSkLT+4a68x9SIpYbt
i6VwJHbn3Fu2DBs+TV3j+M8LgXydEB0a3v/YmC5ps1UhYiqFskbqv9LiVY8t
AE/FBsvc3MJbCwgx/DGUmPfnPNSUQ++Hcb8d8dZAJF5m2NTRtereFH0xsK2+
oESSVeMMBX/ibNYT4D+s3JNXOxha00p50cz+qQeg70FnQvBczor6S8A8f/17
pL6/H5dMOEbKLI3TOKNFfTsQn3L7PhKZlWAUByIoKqL8rDNXlVxJAPyQqSgg
KezHF3J0MjTmHH1sEYXGebfNQ7iYv0VwXeNLJ7WvrPl0B/OvYwSK8nHaB+Em
bayLHSiuAr/ZbXWxxx3mH52dJ5djTJBvNNh8iuwngKq2vqD2TAupD3ygJSDc
hazQv9uu5jpudUjO5rV7xrqWdSQcW89GamzpUK/CPd+KefVu+qJXqX/s8zKv
vNg6B0X/ELmJmjkjdOWgVcIpCnB8M8+8NVb4YTXPUHlH/W41Y3vzqcfcQRKz
syiSmpb0AMlTXEAF17hxcGS0/QsgDca9duLrfmFgvUjbV3d2EQ9RRgy1HzIs
V4pXNs9nkJxDOgAdgCuS/yVuG+OEtLjeLD7mlN94/diTkyznbI93Z8gQgIkV
1RxiILwX30OtVsTu3mPrD/C9CqhlR3ugsd0vI1J1OgNLYP8BasQSerSnK6N9
WN3ogp/g3aQnubfQpj+p8j1VZTH+zAXouLXpnes0Gd7xleCrBFevqRa+KNYM
+3P6NXKtNw2pIDbo/iCkkOEOpOFR3KJ/x9U/43Tp8/V6zhHzi6rnszQs4hip
x9STzgDC36D6P4/cpMyTM74yp8KDHuLCaEf17nFHeyqsgvDKiuzMaW6jgksN
xa9TrV8duLrrUUDlPm19s+wNVVLZezDj88sblRB9LoOUwcChA32QHdYTf023
sgTSSEojMppXQp3V7k4VOAYID0Jww7RfiJgXgZU1v2JGXthzc7i09DVRpm9t
tP7zQeJ1AJYdmjbIa/jBCXfNM38XXcxlRC99EFKAclBifV4z57FU5Vizl/EA
RRIEOXp8o6ScvUJqcFK0PlQVHAT6/0wJiCO4lbCrdgUbV8CiEuRzRygftIst
Gfv6gmNyUHXu+b8cJD6VS2yHZ5Ki0oWpFDGxWNVCpN0C4PlId1vUXFgNObDg
MOXvbvL0BblGn1yDryw07R8DGIU9/pf4ykYFuKeoIpKXiNAqig6D+h0YNZlC
pQQOPxwPPbz4x157wA9sK84FcM0LyNmLsQdwFTbHfMgnyZhfQfPmvgdSojcR
/YAPbuE49EWTRqBO5AL6iGPDjX2NeEOPq6OhNiWpGcrC2mudBoMlO5SAGj7O
VhRoMxi5EilINSGoRNUwyLevdCV0zgP8z9m0tZdO1pvLKbhX5jhQ5NWa4Prf
UWcaahNQovnsStLhxwKTDyUyjzRsmRGFA6DQ2kqBsxiIXQWO8LkqZkGqR/3j
i2rMCkOjzQ6/mGqjffEQrMK/C/lsmuumBugZ2H+irXxVnQ7oY05VO7ojQM0r
B1T46ff6BVK0Ha9sUx2EtM1krNA4E1SP0TWPeO9SWiiYvcltFfNVvD7EHey6
LNgMvvCkkQinoasHO1MSbPfGypXKjCKhoj4BVldms4yktYN9bFSItaiYIKXu
T0ccSXfOapR4FFyZKT4Er1eIMrI7C8bl5BF7JM25enCYqC9lDN3qSeFqOQgb
yiiy6k/vnmjgJA5Q0zdFlw+XrP2MuXIDGIefDvHaw1L+RdVf21EQL9HEVE0v
KCadbHuce0JnMk+Pbc4UMDjoxnA5tgadddP6DqDWGFVjm7v3teYoIIEpHwrc
88RQMz/blfkReAkxJQtB47L4Q+mihkflQpKc6+vlxDKlWs/c6nESLCN/xGQ/
DWEG5eOm1o8ljtNBLunxnB4gyTSK7IvIK/QHvcvT/Cxk1aOPbg+lcHkdpdBg
fLDxnkp3jrvTNCtKB3AU4k/NRn/+QCZHfTRjGsX4OIjeDqTL2TXL6NdNIO0o
NVsIRq6bLOHcNnkWBxrLywJebfkD9c6f9z/gxhhqvvJUrlMJs2jHqKdHNNa2
K1WRA9mEXJcSuIXjhiQEDbLXNfm2jdgHurF8/kg8rAKLjn5WZvoi1JYveeSD
a/LMnygTovo1S0w9hSFuydiA88SzU6PPlX8oTMCRx3NdS+Xl+kaVcDkqPQ+2
CdhOEYCHhL6vF0ok2TffTfkAha1XaH1cz5xB7OKrnRzj/3RRwUZTar/Y5dd1
vIP4CE6RHoQAhqplaZl+JsZOrihkm8nhYzlQIV1CKX5kCxfgwZ1Aqutp1Y2g
yf3sx81GRNyZ/tP4fHA2TME5gIZzef4Oo3U63xwme4qwAD5EwBpRnMsIFoyp
TJI/1jeALiQ7xG0dmcrBDrkvcQDmBbjuyhL34oPCPxY6TyiRSGVqjIq9U6/E
jedM67FEikstN531wwgP3/g4zl+0LMd1T7+3oRokw2F0uf6pe4Rf7uyaRzzD
fOnSasd/Df6jBBCbsaRLqyhBkShdOuMzcEPrhyvirvpBgvLSrhVUacIQ529s
cKSetRG5NRWm4IZTki0lcEWomDuFuCxYKqcvmJjU1PRo0PpVMlUzU2RGCx9L
oY+Rwja16qxOmv+yCOxZqckuutdA3vzjeQNVPCBU+2ILCx0oswf5Aq1OKste
ZZq1SlUI8GjEN7IQN7Q0JyTlvtCcKhyXcgsbQ4Ef56G3VnEtapOL/O+8Jqu5
rogIFFe7g/HVo3WMW0C1F1rKDY1ImPGRldfGIFT5mAx7FNTHMhExJIzn0ObA
dEPIplL7aSBDpCObiB3zEVFpnltryi1iWXdRH9Pq4pA0gWxOHWSLy2NAZU7s
7d+oJWbf+W9tt4fwUfTw74pf5LlvRdzITf47WiFwgpxSdunbpLbeJDiKDJwj
9nWS4oXW+9aoNyFYKn7nOGe0pmFHDYs0hK1XaAfBtyzRED2W0U0EGs5wBXlO
HiG8oCebyPoHPV3+TVK6SuXsLSziN6sFE4E3h+wXexmRAQm2so1S4va7Srcd
LvnSYjVAdNyGKiQmSZc40ylrZD1xuu6m7iOFPEVXJpskUQya9W5Q7mnk0JoU
+VKUzZaGP+aEdGiQT+yM1NeEYOPEAXfiwxdGiKJk+DBM2uHyBmVGvhbYaayp
Xp8AlKbe7SMOm/xrMgVXMl+rZhUqIbT59INtRMFXPMcMTKh3w/Kyu7PXVU/e
9AKHOCHv2Oo3YlVH91ocTAe96Gg2WjxlI97/20GD4s6BAteA60UosrigJCsc
NgNKmc7X+GEkolRnwWeNhIDaDE6q02eHwQLFi2h4qDDDA3HqXL9UPVY60qj6
hkiY1WzWCYbS3AYYAveibTwyaPVTKlNuqytkFh0WbteMB+PZx9U1T1mKzT2x
Eq9ULF2FgtrUyRph2SVEO5skLIpH7j45i9K/+Nz5Th7iv8/UhuS7yCUlOmGT
RNFY1qsf/ND188PssIXMqM4gFp5SZOINBLqt736uay3J1QpWtnxkd93WtBvq
Vr0Zve0Fj/sWy0ZC8CKSo1sgY2FRE+tXYpl9NVeLCsee44O2mD62RXFzwbbw
jG/58M6/8pLx6+1/foVXmPMobS933Sa96fvqZD+w9c1TzhfDsXomfQjeO1Jm
rTZaXgIR3qHCoCePBG2b1/YV7qNRDMY546Ffb7V82BIljJ4IPCueQe1WIubb
pC9xvuhgKke3YW0vIUT8KZx20Vt6sNpMj3mZsjJqe1Q/SOF3Wh/OZOZINwF2
aYNnP9NK+4maD3HLbI5jQD+4ykM+xoRJTCM00Q7hUKnIEwuDHWl52cWIjZZU
2xjsX4iAtpb6TPHGoBoQwHE+JkUttfPjiVXoUxwZzQm20SVbPauhCK31GxIb
9q6U3Lx/e45damrgCbKFMrpFpsOymFAlffC+C4Gtkvba8WA0RH9PHlzcPro0
o7E388ysvsLWvWAPsoEa0WA+OkIKkZGe4gSnCjPep2t036+ksob8stsDNpF2
nErrGpYYiZHzGxfvRv8EaPfFJfEOru1nFIl0U6gsNTppem4JFJDgLoJ16Sh5
NDNOybzeEyUMnEKBVpkftNhHY6RVfZYmUJ8OSTdpvatd3fjF93PN+T0PPPUt
e7RFiE0bhcb7chKdr9dDLjwDEenp8xGavifKMdVkenWCjjtc75IBvVWR7s1z
l2s+Q8s151zy+Ro0N3OV5u8NoA58k7ivrSkn00MbIaWZrWQuOCXyI0PH9M8r
6/bnsEdNi8ECm7Jl+KnwCq5yTWBHGXuE+qKl+OhTSKPUQPcrk6ph+k1aw3ml
6yzuB3h2q1WgYhZvgVUvPkyp8B9ImHRx8psr8oAktGz5ELDRMZDZ39ub2E5E
TgdNsBjxsvVAcEkWhXHGjAsV3iPmKHBhGr4PtU3ZkCxYMJWva6WnHshmCzCE
F5GMRHp1wKXGTuoPnkkMzGLkDS8314n0/xPvDb9ySWFxNVlReboif4jJuoRa
HrF5h5uN4zhE4ZzNR73BMfU1bnrERZ2SERcxVoHz4C4w46IEy3Xzaq1Rd08m
Cpm0SGKmahYTMqGUCwBbRc/EWWze6U/z2MtZ17RMxAt5vvkUX8CYaE1rQiPr
de3ZRGMrxvgjpQzgnkmRsNHgAfGTNRabBo/81CNJYgDXA7luP9YHPXVrCN+o
aecCJwpue7ggoEaW/eAE/SBYnG4VgglTRwA8AehpkXCZb0ULMV2jUmC3mhzz
Sic5lDD+UCMwewFtZ2Lw3/7VHczElnebnmzDW45x16F7x202NkrrDJYS6a32
nutOQLbO3cttTqAFzZ2oI5hcMEuqQc+STArtzR6erCqIcfdTd9L1fz+yPXbD
gHms5oQC9uVxW8ujYKtKLUkZkRkqwUTn9bUYp57ymjK8qKAP15RbKYAnuL/x
zJPLsWlX4Gdu61ymMewIKaMWuUNdjCBZA+gFvh9Gd1TJQWzmvXIULog5f1pT
XL7vOhqLCt05VFvpnda5EpJOjk7FC0TFaFUtKOB1dewLD9Ta8HuQCcg8SYsx
PG4urbnFtInN/DSOKkr/d4fGZRM3eAMtf3EwxAziWhT9mpbSSSd4/8c6rUKv
9L5uu7kFT440Bh7Orl3EzPkWpGHCXIQlwzIVR0ukhTSrxWUlQ9lFTgaE+yiy
GxzU6PJV2he/hFgDHia72by9h16SpfBzczPzSqEEnu0doqUyaKZRJ2PiqJFD
wppZsp/kYtxukjJ5jfMIqyVQKFxRyuBbn21RejsJrWqcYstoO8kKbc2LtRRA
zxXsZeBFgn65LISrM6w1Ejq7wel47RCWcmwKN+OxjL80XEW2+ILkMWjcxau2
cc2qt6zU0byy6sQc1bYeD1u4ypuK0sqAUxnZZyqZTjwU5jVs14PDC6FOAIQf
Qm9gqEPQkcPku+I2BtgIldDpvrLIYhGaT+YAJRP4AZWGdQ7kcFhRlTRkdgmv
ZFYYlAhF2Km3af6qhrsIgCZ1siDcA+9V/EkLcG7u1zHkINWu8jf3t/Jc2Jlr
H5y+hQitKlGhpELq2MLAh7qMqZh+3WMEDSZYyTOjyAIfBEsBiy9Xe5LHjq0x
YbTquo2xxqN/jpN588Ne2YF5mXzhNvxVeRvKzuMTV0F7dqZlLtwGvNi7KdLH
JDBfj++sY6NmceIb6sMuimp6KOSW7UEk7/OOXC54pK1+TssZC1bVhugOaw00
D/EiZmtIHsXRa+C+Odz4BDVOZC4xyaSCMeGt7h+tWT4UIzF3uKi0NSdnuRBR
XygqASYeAKzJpwnXDiWJ6FY1N2Z/SZlR7jjIXLEXw3azzDP4GfV83+g7h5PR
V9ZaPWw4N1Zw+XgxpQutwFEXydXCik5M8tmA+XXqxgb4bUY1M0ZRcKXlQmKP
w1kZtcwHJ5Og6PbgTfN+VvqmmuSsFl3qHiu9m52rVbtvok2YPy6GHqZGApbm
NcIi6tyRyKqNoXwmBAq14LbCWEk+zut97F1HcehXI+y+PbwaVplzc12RRv2G
E42n8Aiby7zqA7CwFENXiDp5cQOPefZyCYp6Mp/RjMpSUiiwkKRwaZ8TIkZv
I6fRjt1YFsSZQkRSpmxCXf6mqpVhmr1MdU4cvmu/Q23FQnl7d+xD5Ytq8OQY
I7oVU7N94kWlppnQYhmDRSRnoPNgcHtXp2w4kjr1LugXhgA3s5LOWj7jrY/C
Er29ts8sr0aMzIP3n0xK8xKPxYS4SQPXur1jXEK9Z24mgjFVSnSBlG4Lpf+a
rVOMFWPOdz+7+IAC3UJ4M2UEk4H7nsnrDuiWCOAiLCntvhoCYBVAvyYkmZZW
HAcTOtnDCihAHpxv99f/4Jqbkg3knPZSyfOVAMnZrnN2HYhk5yttpyuFmHT1
15MWw7vTVXflHvfSRiqJ4TzajhOFBAHA/ztTz2DhQDIFb1w5l/FOcXhMQdex
MWJhfsM9FKDVmjzcDps1rEpdHEc9ca/4NwpPM6x/4oXFC3w6dZRDX4B+BUzY
DAGBOg1RkVmKIHqrbJX3KjNDpCcKDPBI+rzoeXzba/iSnP6qRQ3EIhU/90vm
k92RRTpsPzGzMZdvRAj6Q0TTHAVC+hxWl4wAx3LrvW2l/lcO2bClRC8ECjtB
Hu0NKSIsAt1cXeyHPbC7GeBlitlcYXEMAfHMKipf+U4VD1pMsvaKV6a1H0ZI
H7FuArb8adgZB8FrDsekIdka3eLba8l95q+15TwpZRoX36dE8GbpkxX8jPTC
o3XHtVfDqLEzP4m98qbG8zRVILTNYyvxm25pX085k7pXMBiDRt/hGzoNh8KK
XyEPEyYuWCFEQtrajcCBu6UVK/rnKZ2dPpfqUYU1Jyx9T+BjKWlP6ojP4tvw
aeUsiHlffAIP7EmrPAIkB9CQdoPu2+vuVA2VuA8/vwkZTzR4plEyyipyhDGP
dhJ1QjkO419sCzYFfgXfJfSIjombuwjVfLF2vK0FftPCVk35gEAFrhjjd/ys
J9JleA0g0T4K8VKOZKKHwd+kSrV5E/THPC629eRWSK0sUL8ocxrDgyWEQey4
0FItogpoQ2w4AGYVChcM7XWlOt3cHeamTm2IVN0j5AkFvVsx6abqt8jDCa+9
Pk5KCVYWcCWt8vreKLN0U0CmoXRQyuzmbrGrgTiFkBgfh/8oT9weE8laWq1J
D1aj2uc/UZMHQZIOokC8S2D+GmG3KoDkcXAbYvfhcr3gBFIJRHAVmSUhZNy3
OwTtZhxxIjQd9VanuWdvwD3EIBV+0Eiy4eTs3LhL9W9IkW7zfoK0j+658uu6
uDRxKfYTdzhXyHoU13g4VU/tNvy/t4JzOjCB/xKZrEgyfMu+lEdjXZwmm1vr
Z9IgZxUFNczeZpKi6/4zzlkT48xTpO02rnLG7Ns8XYZLNwChH8PKbPX7+IgZ
u8g5PxyeBKrbOqUGwR/6WX6QsdnFKLGluUyfSHERDeHN8OMECCU+7oThgBiz
diKklA1ygQpDMBXu+pkCASv0O0DJvYFtiCk/OJg0c3/HLIBvYhSXleyFuazF
LDfDAYmd049x0vetnHirxeBiwGbkdgWxiC6istCSQzfT8coIdsyNq0LKw/Xh
MzUs6Ip0VYONkJSkYcO/WJBUyE3Ob5rnasMTZXVgNiBSxPwwNA6r25ql1pTP
VS0jwGT0JHMnj5RXUQUQVV/sbFiEe0EXAWAPgGcIRJ84UO3Cq3xderJ2788M
6MvPPI3lX/DhFwRYn2/2gTCTXzN9o89vY4HTFrff7vUQdSoJwUz9FPJUsVU7
Zc7OEr1TgIHM6l62zUmlLDrI3mqYa0pvGPSSyAhcRPi0Ny2Dr3Hj0IVlVuol
cCEFm5L8ZDZKKTgKbVmQhpSrRXlhJrsuxvs4T9uVIGK9R8pOHMjRohzIfQ2r
DJ0Fnt3IRAX1rgcyJ7ijpOzaZVNNtVhw01XWbSsxSJt9fFqjGWYiddr2e6u6
ul0Z8dat/Dw9gOKMiOMHe01kfxCxjWDSGDhfxCO6cdQW58zPJmgvHLTzRp8c
cRx46htf4HzeWio67/JJ5b+WHKP9eL8Yv6OY5FoHOvqAtRFHURm6PlvQZks9
5RzjeLjObp4IpRRYkb/OoZ4PvHvxCmgpbRN4GF0rbCfshDfV+ffru8DXI03E
Tf7ab0NIUV4HvY15iM/GDAFV7QcrxClFaSUagK24o7ypGGBc26H18jDwfCiV
RRNJ6LRrVa8huvGuORvURJU1LxCF4+Tubzsw0PrlZiuw+gRGIeoYOnwm78/C
Vo4RgFB8eWYpBiQEkv5Wq0MrlNI0U8HwbbJbECJicW5RgD45QIzyoy24oMG/
6NR701NkvDSaeceCc323dYDLY2xrwSAy/GbUkGW+U9iCgd4+VOujtciMrw8t
m1ErwCGamsaopNf2KkpLRw9A0hhI47eNaA4JFX+lcP2RquPYRNnCpjoInlyV
qp0EArxZC0+1BqBOCdcTY1b0thfThTt7vOoQep/4MaR8jhX9cYLjQ2s+PhK6
r+HnYThwryFp3njXEbOwMKtcRXsxFDh99AYSb5ZL6azoVceiRHZifLn1hJEe
fdvxzfQGZb4xvm8GEqaeMbEt6vh9CnqPVpONJFZcWL2O0y+CTYH1F7YwqVro
uiCR6ABheSouQxTe0Hncv/R/WeZmLjTXOK9IjbeDCxd3wK/hplULrkbXe9Ec
9ZLD7DaFhMjLwIJmJZnTC/scBxpSViNmd/J7zjUhJBdgQJwFGTqYGZEHNpuG
0HRKqtMalLwEKKNoq4SEVV0LqCWNnUb0dfKiId27Kepog8AVK2bzO7w1oSoS
cBtlCVPXNkOrKWxJMk5AurSHlogyxFzMel0z1fs+6AHNqRLJIKeVQEQoGFl5
L7XSf7rYBDJvZc6rvHJ71k/FwtHBqFqIJMUva5n7pcPwdI1crANRWUB+4vwC
sxy9sFy7/yW2AQYS6PzHZxovrkXfTkFIJutboNpF4d1keOnvGMXBTW3+tv43
cMYk16CyHM+L0MjPgcebl9Lpx2BcFWZ0Ms0qUoqENWrmAPbMb2HT/N6DKp1e
cHQIZw69SR6AcnkTW1AJpihhVlNsxam6Qackg2+IcuRIiJqMLwvy1e8ggshT
jzkm6Xv/ZPBj2q0+WwCFLvfbty4MowsaWtMDlBj8A0GlS2ac8YERuFQIem1x
lSN/a5wJjaNpXDXfcejgZllb0Ht7B6l8c4dzraYDyeP5K9oM9MmcyZkVXKQV
ZVE/jlbKKIaICJo+HxkwGffMb3zxwKLoIf1yGg8sLMgeL0TH/g3xnwaW/jcR
AQKvglTtFphpfLe0gVFbGwJoJDLx/N2bVBMuIMRqc7e5a9btSEmSjmQCJWhv
DlhKjEE1UJmF0jGctQT/q2S0yak1d6qALzHZVoZHmA12TdQa6nVV6nVXC87c
jJdJLaXS13+SCS0UIKDoRmUXOC5JUGvkbaIcY5ZrppZs28RKUHrdjcVn87sI
OlcaUU85d2NQJEERXzbQltwn+hgyMFxUNOBU7k7C26tv9vtX6+Z7SqliVTkE
nCJoHxU28aNu/9J30Je91V0+FeHrqT2eu0F7z3UEQFAsuOA72fgnU4VK7OH5
37IRIOfrsHzOhzzPNoPPRtn8MqcxCpGTVWX/AzZQo07dXqlx7pbCVSkB8AdH
6Fns6Njm8U4tornT7NecUGNcmHj56/u4Kn/P/1l7pu2nb8A2ReMgQGTMX2vA
224sRklXFcqJ6A7LYoU8/ZRtF0cCqLYe6libOH93aiklt5nqpExf/9tcVR9W
lxnQdkap/2qRzmUv/j46NntHo4J2PxZXQBXJDB0edm0yOVrRpKMc5oC/QQ7O
iZecfpJOR9Upngfy2FYdC2tRksmtGVynpH0lGG3hsKLm1ImMoVzxScMHeLfO
zGTxydZCJtmIe0RcGKwj3PBn2JMnc0ceeop3+yHscQ/WefOq2sg0A9ggu6A7
Xn0PPSPK1cNcTPvT9D1zzHQ++QMnzkYUruABRfIoi04bwC0slUMwPeYLbyqP
DtgKgQKnqfWNZ87tCrWmetopnevNAiPaM4demeR8fqF2I/vuzKztzWKZqgAE
zNJjJ7aqAoAfUkJ/pv9klV7DysCfCceYOLMVzg+iPjyix5lUeH+flgSwF1Mi
X+pSKySNrdZC9kMi0JgLGBlrU37ZxkZIoHmovwU1exLG6TS2cd/krdLfvZOF
VLUsHsSSM3fw85ChpFGzfpeWlPN2yk420CniOvKH/vKIH6dOFRfuassRivmO
nazKKHJpqzupEOlsg8CxIcaZIt7c/7OeQ9BOeBKjIRpD4z2cWgEjMKOuohVl
cz9lZpOYFGqiec3yBVxXbbifXQyrNsq4PuXtvMFNjcKQRwrGIX4KDjA4agoF
F4qMSSB/LO5mtz5Pdy+e/rXb5biYSUq0usvqZeQDP4SJkOGeqiv3Eld/Rue7
+/ETRl4sLitr/vxLWIq0nzTqqfcASb/Ino7P1u1eYtUfs4/3V8kX6fRoC/qj
LJ2L0pyyIt6O/xtWoX7HrAr+Z8B8aLfbJzEFw8NasxkX8bIHJPIJ53+LhP70
C51wyM6YDudL9UpbCo/WMmMi4ZOGqMgn9chuDks7XKUndL2RQcAAgEi1qgVk
3aWDmK88zCwWjDiprZc43g2YLTq7a4q9qOAoknDvJpQhDFIP08HJDCpP2iMA
HcvHgTNX9whXPVp1pyb4j6KrDKdF7i9jeCJqQ8XjkD+Fi3TRA+zzheZcayov
heTndgSNS3xRpGjK5mz/D1BeIeMv4Y4v9OLFRrNwTNBsLjw4pVwYQZyPY3d6
LyghFiKSLRkBFX8/yAyWiBHql4FNmS8kR1Kqy0klI1NqoIRn7OPZ5YidfhS8
1KZZfV9+XC+hCkOKTu0aT3tx5pAOoQ1JzKyhnij55WatbJ+G0CZMW+qDWtdB
pp2Aqx7NXDDrpPLjPCm2pH89+G7wWilx8fldLKy/sJoKWt3z+7X7eAGkmM0L
rqPOibbQXBIOEixRBNRTXvMV+kFCZTNCVXYw3snSFEDSnSf5ec/noNwM/4MQ
S+ducYP+kQLGTG243slJdtDuqgLRYqfnrwq/kv1/5Lq5/wS28QwW0n8fUYkD
EZjGswiKr8+PM4Ep93AFtvr6PJZ/WN+YMx5fK1Y7IgYqsZkGasF23LGDswVh
OoBTZw7YgfzC1sOj3vHBJmSgTObpAZUHbyFFQxNAYbE24gGBVzl/2lgwF/gm
ZqzkDH/pNn6PRVjOvS5mlNmiIKYK46jAg6MD10loRG6Pr+qHUr0dOuSD1bTt
5wGyS4r9Q+Hx8JZ6CghfcejIDzXuQINDlSiHHE61a/+Q54JeVZS/RpoQVNNo
7OF9fS3/Yyfaw3S69TdpYgn0SgziAYa4REPM3leh/AyKtlEv2YyjBh+devyS
1/eDxYOZL68EyLklPBnBwFLoAEpNDcQ9fQAdV5IiG1aVuSpf/EZy+5XLYdqU
5h9NU6H8uk00AJILR6YDnSBCpIfZOVaHQk9STANN99skaZ9Hb+R8O6N9RbQY
rdIJBXlMkV+gMt6HB4pOTYS/pIIA9ELUvNMv9befS3EI7GXe1MXSI8xEeT2n
HtAVZYgAM3YeT9PApQ3DL6ycfwUuM58RuxBZKB9/ISQHlOjXfWsXcppuzFSL
G7J5G99hs+m2ynJMeTguQUf1kOfUH7ximiBZzaLZsVG8vvONX0YqHvDYQfQ8
s5qu6BIl+m1Dc/55izIbLnlhCA1DnWyE/XhvaYKJv2vfMmwlKLPNBd0lWLs2
dd7gAy2WwKzVg+tAJpuf4cCL63xhBUoAeouMMqOKVe9B+jJCWZAzCTXsjGOc
SsMVzHBgIKeQqcpRByWvzk9QvkqJG67G2L2/+YiXRZmAKwcCcTh2O26E/PV7
2GX/9vdWcmBEpmoS7BaLgPFX7QtXU4BN49p4V2DVrRAf68mMn8dxIsCdUoQY
TvdWpNdBHATgMexqpXvjm5dq+sW5BhZc+UMx21Dch9dyASM2Oo0gqmQa8kNU
p9lEBQypmD+UfAYswpsJ0P8taF6caU19o0FeZjW04FO8wzwH/4NHll2sRKqu
TS5A/GOxCVoKVh54jTQSAZ7SoTqu0V2YAOLvw+duH2zcYOozlUN+pNlYIXL8
kHGfNKqqy2lhth1nKwy2jG/RRtvvJeo1wHkF04IIy+sEhETbF8xOqCF4wEbO
4VstQQDjjZpPAbBUji3yrFJhXNsOtF8PJgARMjG34L74z4MWRWhWP5rGdE0T
5Y2TzHpe+SyeUoRkxnjrFXU2iCuffN+tA0zlW+R13t7Gc3W+xgoBOUOaZaXA
+g7YtGFXsh0ciTntsifOK2G1XSVVZOjqGnIpczMjeKTbmd2xW/f4Vqwwp2ub
qgtvmgInmS2Qt8Sqb0Kk1zWnr+/lFBqADt793QvpKJcSed6kCFAHpC9zoXwV
4MlEs0u5GqcmsBkhE3gdoinkIpH15VXID8LupjBpcKon3ckxsX2dl/85O4Tl
BWxlg5Qjct84tP3QFOQ0B/KH5nqqv5tlbhulkgjC2AuCyL/FYFIViZ//2KX5
V0cUfgf+Sh4YSGYonj0EN+4S01jKADRhQpuAZztS2ljH5hjuKIv7nQv2kbwd
8BZCholv5+IyIuRjX28Oky74scY68qK9CPFZIlK1HHj4S3ZQJ6PajjEvUn0P
1FGbD6l70gIIA7GlGwDqLF5e/gQRBf1eWYlkeNWwzvv5v3zZtblFsa/SED5X
fXtEA3Qi25Te2yaUQW6fznWOaRgHywyrvtGpp+wiX49uii3yiXvQwJD87g+t
VqnmIaDmeb0BkxI9fYoE5MLxoXT1YYolgoKlulR9vajGiyo3L6XCU5exW5J4
9ZLeXOekCbNttZM0DAg69BOHVVWFn64d9kOUtHuDCh0p5fc+zP4EtlMsJQNw
CVcfqEUuaoQWLFNggpt0FofeWVsvFQmMJmpfMrw8neNljXAoU+TuDHipQysM
oJsUVV66JoO1/gkXjrCOaADxkCR0+IYIhgi3yIxgnb0eYWwFFl/E1w6vM3T5
J1rkMgdxy5xLaEWKTfF5zSJztKCBf64ynBM7sMq191HGAq4z8CvCoSJbMLDY
QjRUGo0Tb3dMYw7thphl0qQAacalxprsDfQTJmH0xPvHFoHWs+hUNQgW8QEV
9xn4rRb0VveuhKKZDKIwOLW4Dnh0Iwxb4iObv3/zKrESTqUy5NAARY7IY8Y+
LBBfG17gPMMWku6bN9kWSQRDAhEVWSh8y6ijvfuGIDhh7tVTWojryNVYoDsA
wA7mlza/xAQd8enVhYwGa4m5mpKkbFpac+gaNm4bE+CGuBa/2SmdLG6O7cfp
0zK1NmwRabhqmmNcJ9cJYBG4/6nRqFgoMhlaKtoltX9vrlVKXsS+HA+8R+9D
rn7o/bG8CwK15nK+f2koeMKaPSYUpwbcKxDMpgPH1Bnj6hGME1nEgE4nq9Z7
CNiP0P+nmNbijIQIopAASUIABkbmDexo3AA/Io0wxWq2EzrI9N2eO7IB+/cO
1URqGXeYAN2jW2NUmruqe2y+09qBpE6H+SgQ2h/NtbuNIUUBnMES2JB5hv9A
KRhJxj8tZeyc2rdgH+saELTCWpb9j6Kqc6QhhfiQNH7HSIBLM0UQFJvfy7wx
a9j3ADZ03j93vtLI4a/pFEpVXv6k1Lp9Qh8dLq7B3HQt6IgKVVtyapmj8BMb
HJxTv536AV4jKh6ApQCOPwfF5tn96VHp/hGO0q3HGw7hwKIaDJp1INeKk4+M
jD8JkaAagjE38M7qsv+q50r2OSuJGCYRUYpNWw9F5LdAMkMUAVFMTzaKdfJK
FSWr/gpz1EQk6O+hGGQN1rEzs8Xzt9gHzI6UuD37A9CbjIUdhDXwIJjoWGYn
q21TmahXkh+h6XCgu7iMRPEyXuY7/6Cwpn9hyK4cAmnxnE92y9XwmDN+cDBn
pfuqeHuSB605R9VO1pj+MRN2zCWzyWimKLjkamlitGChioPp1KgQ8cxUyGfr
Gdc/C0UhLtOse3EyoKZeyXurJg3zQsN9qTXj5OkT2C8a0rWppqe/Sm8CVqGT
eelMWcBUDExezV9ybDwbZuZOt4/cW5Jsr42zKFgnS38CRCDrKr+Y/+RlHdJt
u1wkz8n2AkGlMoyGvZSFXVRm7Y5JjLVSdPqrPpRC0hcruAi6dxFYn2ttn9g6
pxPu6Au9wk5137GMGYcpONHpxgMeIcRkizTFZavd9dosybdPSGxY6AHnniXX
3EdEYU9ynWJpTCy4as68lVeDaZcYcdyCu026tq283bxxYo84XvC9pf18OcHt
gNBlzWFdKOR/EYMvE1rOrIsATuPtjjYtYrigPPjcRd0DMrycc16z1vT2WyCL
iEs+ndjr2ytg5DNisRlmeFZ5HeRH9IRPeFj3YyzqevbxhDDn41Mp4UCzBhbv
KM9XF2gkbXoftKAL1oQa6vqItmvkn1Ner/+BrAS1k7gcINEUr6AN8PSeRYxq
RzIEkhxpNkM/SQm0DOdMOT8hOyWt8DnhUn4qnoIrh+fUZA3r1rOqJL2yuWyB
4oMvN6R7bSNP+pwQ45G4+6NJI7OL8e3dSohLzs4Q5yj2lnzVc8mgXRieNxrH
3QzfDT9lh0DG1qmuo9Y/0Qh0j+HbpYknl66fuUoarfb1h6fpsQT3ckR+7tCc
RR6kMS2H5qAPCTxVD4Ipz2MVmOXNjLml5qPAfpEtkf1J9kuLDN9hdpKa0bV1
JZP9pqU9v5qY9AExQE9K+iJnZ3nRJSEOReUczzPPDSo/8Auj9Zar2AeWPjrE
gRsST0B/XIHf84MxrwcbcmYrVaVAhnbFojZufJsrUExHhxFRHeiK84e8mnbG
gN6SUFD9b41eB8P+1f/TfMjrHs3heQd1TVjg6Kuhl6hIruAG42JgxZLdf2/h
11zgKRmCHPjW9cch3cipDGAKaqUitGekCh8mATlkCn29FzdZda5ipoEtSV2U
l1MPLaY8zD9hikS+ImyDW/BKexR9Q5B56Cm2H8qffY1p9zz84qBphQh9x9LF
yCorig8uLysmkjexsjI7g2+U7wpSixfP1iifRVl5RAtrSLimZ+5U4QeQ2XNH
FThm7dWWi56gjQVIYoTpD+HAJzKBB71ewtkrizCdsyWHRO42jxdpeMjlXXbE
R9QqQs5UEaio5qGAERJSmZHU29Jq4x+GViTJ24SHG5AHi3rkYMP1bB11bWRc
IhyxSr53iSYY7smF3VyBvHOWWw8emRLMBjBYjSKYJkDPnxIicAb4fn/j0VJv
DZ4eLRa4+ZSs4+hGio41XWMKagDnVWHjqI3AqwUesESrNA3ELyOGe8zYLYIF
pgAArlNPkXO6WIFZmU+TsTo9/XEEBhqT6i/boyOM0XE8HSxEb+2hi93jw9Ec
9JDIev5rQKV6JZ2zAOkxSYgI7JCv7nUZRuWC24jYghETZO+8LlPBQw2oGRkW
Quinv8oqgFV519DrfLZwUlNwL9WtmsDYOkSiOJ5zTL6mc7DiNxc9kRxIIH27
AxEMynNcBhVDWpc5BMFTKGOz80ChGz3CjCUcBJCTmDyg0BDA2ebJ9YxYJbFM
HQFhamn76H6XTzYbfSa7+5a6QpcFEpDjANvND2qp69+4lbuLfokJ38BGjC4d
m7WTjZe4Cqs4QWaDEAiWy8aD0ef7w37uAlRsM63P3ZiWSj50KRBGMNdBcPLn
cc+heZP/UDymp7+wdCzhONP3GKB+zEfSyNDF4vH1HUpOwu0kRFj7q7cxm8Vy
vfed0oEG354jPhJP7+CLtpVa8d5Xo1FKhudIgP7Uc1FU5I/7+tFfaaYaRMIr
B4CseevnmvD2kCaDJg0BaCCxc2y/H9k0vzAW86os+09VeYB6yiBbrMufZPC+
YVOf0zSvfwL50qCy1WNWAXh0se4mbUf2ctriHLKuWZ13O/GWThkpTLHSyvlk
K7uT7fQvVBNcB7m0pWQ5VrxFBMAzgnCGy0ijvsMc9b70IlH48seaSioF/fJ6
8eneGh+rFfxjBQQOhCv5fYT87+xeD38KQHppqCLQehuU5IujzKPTmy0gAxX9
B1ijXTksuuTciIkv0/47QJOGmoYbrSv0dlDF7vcYVhSNmoFkOmTx2s3b9xlG
leW58N14mDDraCMxdocU76NOWUaq3fPS9vtNTG0Q0HzL9ikjPHb2HrXqKQCi
myrOEOmnFrJ3WhlO3TthXqn9uYLNJdslLZCC2p050oKvavVzTzGXXcKD4ZNc
QtMa17mVDdKATH71RgbipnoifPzSAnvAd3qxndBBmbwJIT0M1fpcYlqQJ0TE
1dI8ve5jVQylBHaBzViAGyttFc1qGDdBfi0p08hFFLrA55p/T6DdPTR4R6Fy
WHb2i+lVAOMyYqgjIKUjeGhjeze/gVrd+1uy3SSlNE6EUDY8zGXcIj55POmu
jFIo6biJ9pzF+LXx4eyFv5ppLXr3co9DBqPHAqIE675dD6QzHt0rDWtXsMpU
3tGmY7GhKhaNJjC4bPVTW1WyIFdA2KBZO8HYi65sbpa1LrkZvoN0k/d8d268
i0hpg5q6eFtbyNajBMRBSrumbjQX3etGZOBzsX5V+GNMDUqlHZEkv3xmh6EQ
1h3N/v0fqukwlUZOi6pk4KnmT4aCgLpi1B5Nv2VVJ21I1BTGDysn4Ppz0EL5
pmxWbMszng3AdYx10/xAk2B4YpyVpNSZULVtwtkGPmGejRtytRzZShkqKp7V
jNxs8m7GZUED4rfWIWx1PaoyPFN19ej0aein1ZPMPLQmbWjEvIKul7ZTpFoN
13dgU2rZgA1Mjp/TEiJDT6KxLyFXAxZ/JWkgc9OjHMmoZDxFMPKJwcUhSmL9
bJj/MPtIkWXknnEOk9GfA5OvXRfuxn0WSsqogsz2WHdOGjozX1/1YeMlbaC7
p8LoUkcgES543OwNw1FUIkXGBvKEBZFUp+ms4Pltygr/5FC32ZnlVcrw6O3p
/Tu6pYu64S+5koDUH5a3vNEiWjeROi6xjaNLvbAsGJW2VtJKlzZ4r2+Gih/v
cMcOLcWWdLNLDH9b1cAYWumZoVqEOwVQ6KS/NeGdp2InidcvS+o8lEl1XkHh
ibJfqwg33TzMe21i3+2LICdJPrSqZ/v1u0xwBsJZd17UveztWlMdnU1WsmzU
SJNyKxGIa+hR7ehUCW4jj4lGPPHLR9gsm+JTiFD0+QhPJn5Uvhlqg3sWJUOb
fHvbD0YUuAmpSNL2s5P/oseAsajlEd34gDUoJTPMOn+68oCk0LrX0fuygg4o
pQAbHs9LdYGZ/zoBDkYlzRURPVINb+1Mt4KE4ovbVyPdOHHPvMjbZL+3VnRy
7gTBVSMJF1bfJ5DNaae/CLdmFNA7lLM/f9bw8oIZ2wUUr/9/sIKzciry2nsc
s/cKIsDP6FDIYqK2tX2PV0WO/ffrgDOSybLY4fCaLaJGycap5hDbbBOq8Ca9
MS57tFBlLphHDDiiNgYEfAKtKjMXCUFVJY7ZTAyeFrHqyIVL89hqndc49yeN
a1PD7vzjA28O4Yl/GbzigXDFXr4k1N/SyBDCqxkv7/vb3xTIDnDZ4UO7IN69
U+TNojmKhukDIpA1NpXjuTsD65bfFpki+FSMRdu/wFcfOVmq+F/fN7S9gKSe
pBpr7qUEOUpcZd8dVxEsxUgxI1eQ8MzIJIQJ20HH7hCe2h9jop2AefHAEbRt
f49fkiqECy9sFcibqsGZUHzVKVK4JpA45ztpQzafGCCEghu+jZlXHHDhMkZa
1NC40oLDlRPr8fwGhfH3BHgvu5+2Sj5mCiH0eVuz6yotjmC6xc9qEvIseXDy
uSPfJFkh1PR2vg4eL+DlYxbqZyJgkjDYprp1jtAYpSctdFXu/vbtS6hMMr8u
upmNy2dSQT8HNjoI6K5BGcLQID62G7HOoEVJ4paKexVgTzTDkFHHOXcl8D2r
8NLRBy2ZqjMbzgmKcUZZ5y7ic7gGRlxQNbDFVlWHpLiVCf5HMxEB7lhBBtTi
nSQtwHV/I8+WfcuSKPzZR+BT7lDCkx8xbS+U0mBtDLPlkzlhGaCnc/wpM2fE
DdPDCd75tUY+h+lpMRll+8sGiNb9MPGwkm/nBEYElo6jbcPL8ROqYGerkwQT
zVy2OoWLb0yb27EC54osHjBryp3T1kZXxTY9OOAJmtKUsbeIefsNY9R2tl6x
acsdmNtfmZZ3xvVqs0fe9h/cV3Q4gSvJ16IS23f0YQBCSeyCKkXqCQ43N6y2
ScrnAY5tThM0d1gHcMGGwm/Fr64CY8JY1V5k/lNrVVfSE/XLUijrqP3yaHY9
7g/T25i3nAtx88teqsnn0JHOQesGY++AChb9N3mS3SXBO1RAsztVQUSQpZ6N
Cj6KMywzsSOIb6jNrRVD80PHazlrcC7sv2qwAIrRUvHWeEChBkAjYPHVLePy
XJjzFJDf6/SUY6Kc/n9u+/BjP9fCHvr6BkjauOH0KjNHH7c+AcC8F7YPLn+J
eSVJVgC2qHbvjEUOT0p4SQaiM6ZIx24IaB6493TrcJ2JoXgZYmoVAjuvvaWe
ym6qq/vkqIciZM8Y+7xRejlXPXEvdnkppfGN1xmnqEHJdsQyVSt8vLh4jrhS
EKUfF3OZ7g/uA7YoUDhdUonCvldl/TDcSJWPRn3iu7QMCV2Fb2WQ1SNCqFtc
l5vgvGlGO9pUUTjCRUjuhcYUXxLUIDdkLnPU2qHwi7ms/zxcSiWZ2SXwHU2y
r5AF0rAsZc1S+C0jw39C6sPGwdUuobkRboD7A6qJg2KHmtc7UosS4byAlkX8
yFJh7yPkbONytgpgn666XaWXRLJyfM76SQfgmU39otudsq3Poj8FORubgSmz
sFI61m0GJuZTjdt8zjUTzo8JzSCfbKvahhEbSlMrF072gGLGYLVvIT9JQ6jo
AiVXybgU/uv0b2dEmbBKemyhsav3pP8fUY0zfLS0uOB0IR59NXW3k+JaJsZL
76ciuIXi9YpgxqPHwwyjLkmo6wPjU00rZUpVK+nAYHE/OOTGCQX7faaQquZA
YdGbvqa79mBl0ohQZzT+RJ7i6b+Z2Zz4LeYZ4akT/l9Z5OGD7F/4vJxpX0NN
C+nfaX+yr8JL5zApolbYAzS69Cd6omQRKMi+bn17SKvhehjqtb5wWFwyqkDs
3H6buMi0lvt4CT6JZy5XWt3NiCmyAgddLWHbJt0rD+KCvEz7FuQUryzjarcH
vd+ywOmJEwRW9ISySdhrtqALMKsQJigii9iaCXfa5CJA5atqXC6lYFF/vubv
9F6QT4tW/54Vhnfl12KeqUFeA5KKOt5Hjrj0LNYRdv7KEV/6tSgSKtyPdcqS
wTnO3TrFore5d84q2ZjiWoQKZ8qKCgeIgTp72hP56DUCFNifWICaKE3cB+PE
478nmyYP0lIzQs2riFodEcQDyJN14p3+YfkUlyb4e1hSU41RKoPLf11u9vRG
nK9P/gzbgOEAmom3haQS9v/Lor62e6SJwH3KRFRdfbuBPjw7U4Pr0nXfXNLv
pCCuQ6luAkabBrmzREzdp02oOWQxNn1dNKQrUYHofq45aNRqd+hPXJaSkq46
+PbWBrqz1RGhs8gEorM0zxRt7q2UglekW7MIHhKyVc/ztG9vOlOj8e/fGRSt
zKqFR6mPNKtx9fsECMkrm+sCoDgMllv1mpm45jrd0uYfkB3jPItVti7ezTyn
Y769wrCqmg2DFgzKnB9xl7nPFagHDx/Fp2cYq/5/bNef9r0hCuygCH5oWFGe
/kfWB1D2LkWjPiXKrZLOv9s4tew/SOB7zxq6p1FIhV/A6MvLwPUYBFU9hk4Z
Qy7wZ16YGVU9btv80IM6F1qtWHFvf8HnrU24tiUBWzFw/edPvbhcDzHtiTyk
/agNXeolxqFYVqNPOWCj8SyTbPFSBOPjFr8qjyGclI3GZR2MyvL7Vv7MIotN
b3TVOxF5qGGsHZDHNv1JBNtGK2quRC0DbEs9rhjMzU5VXkWErpdBlxK+el7h
+KwPt1I6eDpUFtxm+YayxYNiNhKbrvwHWNsPkewLRbcQ2edjXIGZYmG42WKz
l51xBZDnfePeC6CJ87WydEqb6FKI46QuXQiM36d0c+AaeUqPCdnzd3hO2STv
h2t18laY1Hr+kRrEruWB/i4tupDKnf3eldoAAKhCorAzj+DhH3PwTo06L5jg
1kakXt+7aM0QSITtCGT5pcIKgC+sEeFh7YP53mIUjKFyHr/5Pq1bBF4s/53l
+pIFNTxsYeSD24UndzbzB8djHEob2gvnsmu/YJVH3TUyc1SelYrv5l64oYmz
SqGH24eCHAUQgqtpfN+0b0r07JPzhmIR7goqeA9B+h5iS1iYQVstWLr6yrnR
jF9+woladJcUp16mK9At55zOsosmPI8Q4j+czgJtCXrfp89wfLJt01kApuHn
b34hXpNg8u1M/RmxQ6426uHawD0OWO1dsbdzpYXsxqWxG/HTt6HGyChdGzwo
+h9cMJ/79iSaqXIOBtehaTZsf9/U9kxeEJFkmwg3A+QHrmnm27joscZN41yw
NQiTUoDk0tJG5fr7ZMY7ZbI+tlnfqR5dm/599LJt8nhmrKqfsGSQKwlh8P89
9AbTGDSu6619qG7clBuTP0Ti1GwHFkAKClYIAOD8Dux3rwn3+29mMz1BrBdK
y2Mkz30ra+Daj7YzA7xDeOvNhzn4sCihw6SagbrmDDQCsbZEIUvwOKABN5hL
6RK5VSwc98N0cSzxYIihD0bgXFimPRN2ds5GJ7x/kvBFz10Uz5Pkz1LE9mKi
Nbez27eAAvHFSWk6VYkZMaT6/Z81ER8VKi1m0d7nLlbJaFxmXuv6dmtnwB/J
16l/Ck+hJibO3MybdorgDEXd3R6paARRtriLx3oA/F1YZyxY3X+k4SEEkw/v
/Lc7EzYIU6GM/aHPTr0D8tuVk6LtsA9EyPPz68V7AAorE8/korKBwz7yYrI1
jWWyCBD88goRDpeeB0D9KdOMEWRVpO6kq7JtWgGj6unkgd4TMg5Vt7qoQkR6
8kx8OsTBNj0J2AcZd8IwtwfYeYZzoSBQVk8yuaRmb5luo1mZrYq9l3nzsRad
4i2lDfy0VRrDFd1qW0OmFfe9XNfnyfwMThvtNUQd4trJmQLpRDS25CgYIRS0
ldJXK908GhEoPy0wgPJvIgAo+ALCs108Vlu+25eW+h4esTj0oZ9bVZ4avGGa
aTOe9P/NpVIVlnGeshrmP3SvrWrWX6jUYKYgYJBT3tk6w8jTjUikhGmz+9I9
F0W7rzGFVFIcvaU8/rUszWeZ1lN9WOdvZMrxqlbVYM5qJuSua5dkGPvscQnZ
yj3CKLC7UXadm7GVnrvHcqY1ZSVne0Aq8pcKaLj+StPgRd6rNxH7hrBkCinn
zLuvSNMLwCWWqV2e33Pi2fkmPVLSShDWxEzqnwhDZQSfOlAw0ZgBxfP2oaPy
rwfW17epcS1T3N8VisIgkQo2YAzDP/ar5r0hJ8gByamDFTDcCdECUyhdJZX1
F+Li39RxJOANPXY95QKZTkyU+AVqt8PfHFCAd4N1z3G3n053bHNsyTt9k+69
wZSMWtIYc07Y+rXXRW9+SOm3ywW3kRAkoRjaeJUQazVYiC0uHsqKk2kcke9S
MG0Z+y7Tu03w7weguSy/C3YOjM6BgjkBDSaAwA8IhszJ7tTPosjhlNKYayzI
Linkw74VRpzQV8KhQCQhDJcz+pALwKq5CWRhag8AGCOnPZ1umo1tHUc4vmdQ
brU5otDVaRT2Z8+KhFZqkUZChxRhFlmadpYYs99kih0YhdnKZtJeyPlrRcZ5
ppDUHaa94SzelKE7urfolk7fFdfgAqRFS5HITKD4+zxqSFMZccYB6f2MOeU8
V9EzRzFiwQ4/7FUXUajdLVFkbmzZ2i5AVqr3Wen2x+Wxmzq/Nx8Euxs4rgTQ
Yz/KThSWbcLwZ8qEHfyX5rX/i0jn51kS6MngzuEM82P6+IZ5AoXTxPwXU1+1
ngkzimMMds6ornGIkQHY8lSOPAklEOJGXWAzTmBg9UK6e9Sy1F0CLtofgGZd
ixzPqR3TBOhALfvba/T8EGLGNH/jRv5lEqfdPRvnjI5zden5zL7/8L9NYr5h
eHJ+wNu3UWaWR/Kyt+RykX8p3BfZ/v1CZVASmpt/+eMZe0/GC4hk+/AYIOCo
6H9/I4kiw03CbeiX3QRT1KxlBDDSWAgv1QStPzy88m8Go0xqa3XCGf4QBMnF
wP1UDOP0OAPRAQX90YeLJRymi4kkiV/jxfHsnOBQQ0UGqW9JyYTKgouT3pcy
d3bJaongshKCu9Lz6+p0pO84DKKIrr7p6xuAWwYCcyLawCY2B4ZxEavvECpv
9W8vinxVVPtz/lQtCLP2NeKYLdzI2HV4GOSHv917vZET58m3+sHgvb8oQTm2
Vy5LAEC9RB8lL/+pCgrHLiqNQ+WLL40jpq66h1iGFo0io8yXAzsILBFCq7De
vHKkZf5slyO0kaATTdUzaJuSdzlOxU8oG6ULs8H/PjIybG8jjHKMXzC0IG5s
NnlOnmrk709urMxnQ6Cx90aGmqu2H703568HUyNMbx/WBHiNHL3cdsBQ0eob
wIpXEqYyDtmPuh0siSm0VjoR/rpGZ54ItptTIugSvVMNjBIpoM+sQ++Oe1yb
bOiqkqrTshYIKtHHj4tvxCqK6kO9B+2o9qs3EJ5Sp27Z0tEjCNK5Wt6+g2KH
lLs+UKgBD6OszvWVZRaIv3Zk3JSP32xoJRpOtPiK65XHgCQ+qIWM040EFiaQ
DfzijQcwLf0EQLY2VBR2icm+QTv1aQJ6DBeglJtCjxuKbkuUjNbmxrScwtyU
0ABGCeETncIO+vITHD7y/CTQtWH6/AeNt5a432TBCzZ4KcUOBrL9DCZbVhpa
6N4UMpArP+BbqkxKglKx31z+E1Ub5QHR9oQOIE417I48FXCNCnIxew5KD4Gk
xmaAPFeOUUcPo+wruUqFfpdegRwq8GtxmknrsxeOZBSlTy7wLLOE58R6yGnF
gVOIey3FeG8FT9T6spAJBbRU/Uxf5QGbXsk8NkdXCY1+ORm8deJuw2td+IUL
I+71A5OSCTJboA0uCQnPorpcCsrsqrI+T7imyLibe9B4yJiPYNwPwDTWwa3T
npVmv+cObQnR7d6PjNs7juTGK5IKOAM/Dwt8nhTTzqng5x2E1r79Hp0i3D7U
a3oviONYXySwl2o0JV1DSb4xomwt+UpsFSJZMk6w/tqhVFFdGTzpQOuXYaOJ
yNQigJchFCUmr1jNyVDARe+D4cdZy0pahDjp08Qm/frR3a3SrbLOOsG13GPH
R+ZPj06JsCBI1NmNs4AcXzdvfn/KzJ/g3+Zy3RvjLSHZPGb4wnNbuOwAQ/2j
vosGWYD+M9zQ26rw7MnrBaHDtcre0gT9rAhubToG7t+LZkjpPVF48e31nn5v
aCFDCzIhJqY6yLN2FfPPzQ4BzVZmnm9yofpelW5H4Ny6vocq2XI8f7siuqEV
WF/F6zFmsNoVWrl3ayGsJE9myGApvLdfNn32j8sS/rLUT3dkoYYFN/w2UfmU
lWsyFtl//JxH/PxLz5q8/b3rVu8eoH+aQ8FHKzYMgyVWQR20okZLBgupXsmr
9zD+XS5GT3cj8Rm+qtm+sOhWKLY0KOS0wwlCXbSttog8MRlUDj1ROZBe8zL1
C+cq0oKjiLK7DGGBLtxnW/ywTGKlkoO0twKwGKtjBdPKO2rVXLpSXs+TXxJj
ZbHQ6ZhsvJU+W8792r2Gh/y3tZ073y4vzGHHHSl0s7Vv9TbhDOwxNyqRa0nG
9+pFwzfY7Rl3b9iznfe2J51BXxLalNc45CXxXnVhXvjkJeWEBjkYgR7O1o2N
ZRVWdndFR0VLkNluweELkU5qxhyUkOJg+Y90WQ9s6Xj0CyAQtAxJyxvkDV3O
ZxSmXy6pH4jcLF+HTLDLF2GQgxTTkU798FdvyXJATnYS89/RnokzuBPoFDQv
2yaujM9JU0x01+i+iJEIeYtc/+FRIK19wy6hj8CB+OcftCfowmWi+vJgLJOf
yp4zcImfQfnXpFpCsdPf0+X8ISqFFBiUBJdov8CL6h5yYGvQOyX/qiOGR0Nq
EGkRNHDWQnBpD8S3wT7nHoKsb+1OFAZqqfeg5vNoABjmTF9sv9B3OXO4ePtk
JOvdHq5Oh/+0bTaUj9Z/L9M5y+ZFkQblENO95cvexvmEPXCRP26xdmqwSvSj
kVbHTIMrwyNtNOoXpq9PPMe/FTX4R0OET1IgFV6684Jq/ktEQQH41h8iblt9
s43bnM/hWe6JXAmpJhZFKeC+IWHxQJBNMudBr2P0ODBk2nlKhVzdrLdC4sSr
JvTZTMCP5XvlUZNGm8Cez0EjqZRViFBEprYtZvYQoFwa8GVJkypLyQ4OlQCf
K9jPTHMfHZ9zEUDJf71LQB9lUNhW5mx4OelxdvkF0BM/jDOWQorVY3SF89aN
CaIY9yfn3q3BzVaJPeulDtvQM9HloJkCAvNaVP+vlp5hk+tXx9DCiRiJHGKD
TVtK9xIz/sFrHr7cxIl2f5E7Tnnw+tMD2Apb/FCAO5+Pj9xSNHSk6m4ESxyp
efuEpX7pS4wjs0n0rx0G0AJgPZf/uqcMjLEdMIgKO7q3FX1Y4yh983cBMNBB
R5u8skYlr821OjNDlY4LnInJeyiFFuvoshi26j5bAKaGzsQKvuC7UpDDKOfb
uxnSVPZGZfmGmrI8LDhntNMp3u6dNmTSgvCja2457slkk5aIMy+iB3zIj0CF
GAQSpKPRH+mKv+PkEXHJVefL1ecy4xYH+ElakTm/XGlg83UgYGCLzJWjpBhw
gQ1UN6bqVGu00mFVcuMMd/sd7sfQ+5tbM0MMsZzE7a9FcR/ILU/u0srU0Hvl
aFBEkUh3eJlWDYzGKNj1mYrtM6qC+FLzuTXZcB9kwOYzygRmOpRUB3OYbQOm
8vbtfWTEd/hM8xqHq56Yvr5MgbWDc9WMoGqO3gURysxaQClNPcmbCTLuk4ro
OJn/6ks+ZrG90EeGfYeS9cjaHI/o5DRZ89SrxD4T2l56QZLx6013UKPVrI1m
p85yAoUZxP3KKQZSTEsEwpM0UgYrTtJxw/0YX+HwLLJna472LGm42SRA3f3g
MEG68o4YgLdqW5j9Me/m7lK3D2tqMz7mILwM9x2doVMqfLP0JVoxv72s7m4X
espANg9DBQzRhDkel56fVKdq/iJR+ugQgcN0CfR2xOKs33TNvpqfbys+Ety3
9ju9oCAGQ3wfPBV/scW45+umQByZmGilrn7pRKJm1+LFYhxjgJ689bwRAVEa
ohv4AT7CESrZkOGSUfaoimfV5eGiRYct/ruGo6kB6q8jTRWbzvXz+54MAwpo
d6GMY9HLp5Sqc+aTqQ//h2kDb4IZ9h6P0fSnj0TYqYrHO1UzMg4vhi89iQKz
fbeXZt0YWbu6S4wyihFQwpk+by38tivLBiuvVLxQS6LgtR3bKEIDQB981YXV
p7GF6im3myXPl1lHgGBwiLT1PkudDoaMagyfLy0DMcJk4V621LuZP4Vox6nK
XS6j+xD+GQCf0hDuHletE/fIU1lErXWCqIqW2FgOj7ZPo52JWkmlXRtxGYRH
UAOA8tokBscWvW8szAaYNCBPgv/aEkqXrLvvrgkwywW+QSbIHfO7jVvqXkIN
RtXQBFAc1bzqpHWff5TbG9XFUzQ8BTcfYj/aikpmbrzVw3kOoEKMdzBkGS/Z
e4gHiL/gfXBHjLFjbdc4PRigAYbHCLUSepzh/gmTzGn/4zaO4m8mRFAW2zQ1
hT5HZuDctQ1XRBCPdAaybsh7ObK4X/bIE8XRTlZIKsLEhESuPtr1pA6rDO2c
eghiMDu183ehy9ZkPS1LUtB5WPXtdt3p4vvnLvaJlD4A3Q86t7O9oa/WurHN
vic046Mz1CdaEs3+d9pIylRoJB3w2wW52DFn0kykhz1sHb7Bf5i88Hn6LS5a
Cw6lDpEHvhxN4R7GeI4CA2JWknCuJqe4rhwV2RK56CxwUXcWhSi31Gb9RUeC
FgBlswTFOtPFNwltfp9BmBY/tSLbRIW4M4l5J5zBbp9rM69zuGNRnsV7cnnm
0Oa8DLn/vbDpSDqbbpbFv6b0okEpZxIn6tLgneyruX8vvwHngieAYnoBv0Hq
MmhVU6U58Ga5gYDKx5mg8dOPSXFTjQwHxvwDSFaMYbgl7Eise5TwOO1gMU4f
nrN7x2DQt1Ey5CLOL7irHsNfKpHckwLGTMhhDSpK47AuZv3MBUMjs7VDGPjG
iMyjYvM9zbmDn0jxoO4XCoUpdVocGNHUY5/DGaW0ah9TbYwDMP/TSPgSnxq1
WMxkgYcEZNDUpyJg3VK+8avgnJ2NuPxEOLoKqdYOfUlODnqaATojSOL945qn
tGMnHaFRn1WfJdoX5m7QB/uk5k6/WZC9LAIhLUNhDc30oShgFjBKXhQ1WyVN
AP7Ow1++nYlDOfUohMDDwxsuG0akqX0EYeWyR9znfPIo9jF0Od4ITVw2Z+D+
ltOvWLAmCGDn+O/84h7dR+bJbBmuW4tGqryHBAReuyImn1C5/8djyIAI/IMu
o+a2HsBzeyPqhSrdPfQAnF9TH0zusWkJTkg+AkNzKHo7madYOz+Z+OZkdyhA
CJXOVQTXTwHQQBzPkoRznkccCOs91xc7gT16AcY0Qgngto5Cml0PQv2PXMhU
vaDAOfCjfUcwZ2RknNLSRfBsrAmwt0pQsrJYtuHpiNQYQ53hztiMnxfCVbDH
MQACyjdP3FO0d8njc8JiPBpvf3dwWtm5bAc8MgM7kUVA0NluNDIpf7Ya0bDY
o3GBsMEc0IJg/2kzQwI/sz6AtYqpvpYuRRL1RyBfSKsXTTzAa03aOzWvkx5k
dF086LHtJ9RJ+ecoLj0goTNn/AJQwXLk6oyBgf1mQzYX1qEy8uWjp6wVZk/k
r5qTsnbHrkYAWUJR/3fX05OmY7eu7aDrQ6G4K6GuP/XPrlRDaPHwt/ooi1dH
zw/9mxFDNlX4OP4OHx9O/KM7YoPA6u560trWf+sffasVnVwRDq5qGi+GVNQB
i6J8EsdpuYwx8fKJFEB9jF3JOd7La8pSE2UFfdRqva61QoJ6y2pmoegw2n1B
xll2qksxwfvfye11yATbEUuAaxnDzsQtEMXYcjUDq7wNyX6mnWk8aWLU9Glw
aevy+VwzFRTZjP20GUwd/gV7s36WlKMNcp4iBMC/6zXESVETPo3MpoGl2rE8
ap5aw/5HKPMU8JiLRxOR+uGlS7YDZ29fMru4q8I/niHhPSpK4YBOaV5KsaEt
t+Xk9g9SqnAEF1kAxF/s/c75MTPBEC5PT6DS7aI5iCC1CCQhR/G72zFq5SyC
COGd4BZ4Jm8iFwm5ZgS7D45ncTJXOvWGWw8prjQgf4heZQcVv92tWsLSxYAM
1vM6jUM8HEU1taWhPYwi+L7gCpJTgogk/NEhPrZoAgJjjr1g73Rfjeq0sQZT
hbdPj7RBKCxzlaza/ZhqSLphZSL1aNQbLOvh4Y2bjvqhbR+UByJkGKlDMl8b
Mvega/GQrvyvcm1eO2JfVC4xtdjqpMWyYQ+avDv44LMYgStPEOpR3GIFcr63
RQFIoSX6LgURTu7KF1EHFWKeymN0e6uSkQNdKmfv7nSO7b155NwcEYbaWzhl
lOoxGpeDAYSClXy4cgdKmVxwXBs8/Z1BNmPXQvIDcFsjzLnZjlSQQfQuFPO7
fTi/5fJ3Qfsf/Oc5+DBvVTAuiWkiEPpOYVpOJsecunyFfoH0qf7/36qnSNSX
JsmsV2uubyQJJmfTnz4I/QUZMRj5vRa1QPRovGTmo7AaqL731T9JXPTAKrEK
AJ3Hk1oqTbq4riyY6cp7UkT2vLKgdpzcBDx+QMT82lkernl7R0OACNJtAWEC
qRNDn3MYOh0VxqtNi30GqxH+YoqYBfBlD3NoW2sh7yTkxXwh47C5qy85M4BR
pb8CaEAjmcGe8gRtAIu8DOZHwlur5AWrDOeiiaKdbMZE94e+IW5ndcxcvXLu
XZdzLP4OVf2zqbRIlY7Epy6cwmdzrUNy4yBlx63GWx8ZfuqjhJB6bPvXwzYA
QPfx3Rb8soqhbVPokpT/FnBilpwrFoFopKoIAutOK7SonjSMRlYDxJZdCtfX
TljdxNXXKK1KdP0AfRRS7+1TCZGkaCi8qzc4vMeIiWLZwCKmA6giOxFSR8fW
9nDXjGAnIgSedLTl+96OWfx3MyVXK+o8DbmRJDuCxsTA2IGhC6VqmvBsIHkF
nIouFaOqxQsXH7y2Fp6wWRCDkyPnOEdS7w5PfgAjV/4n2S3Cqe2OaA6dUnOj
tEH1AgI27ZAbtxhGLSHG1YTj6hmoSkJz9G6HKRzRjNWHv/8Z+PRw+r97f3RV
Sq2+aY4Nhdh/jUQG4bEoFkhebQheMmpDZCSvbHyrL1iqt6JnkyYguiRnJ2yG
9ExFKUUB5huj64EDvsiZUNTf4AnB4IAT1YiT8IgXFfYT5GnYlgMgGeGarNhK
0m+CzA8JqIoqLCQDt5MHORKJevwFvtZGc1Qy+DnPhcZ3UooM/C7ZqUiCG+Mb
9/GthDityquR3xJPzvhCZ6OFPjCp5yafxUchFCK87bF0WgfLlZDvmkNbTQLM
gizDvmPNVoKdUwShckfHDGI0vmyMU0MzGd7lVq7jXpWqDLxvjMQwomG+IcWq
XCviyhDwl5L2liXnM6sjnbkqmAMrpAnabryDlBev61A0JbgReqGyL/ksm3H7
qEUI6OUVpLYDF/Gciheax1zAxI2RWh2wDRZj7mTc5zxGic3qhEk3f4FerZus
soSrVQPIyKmef10XfP8ZvQ6gsukPZNYu7SvqyCKxE8oQzA/yHMTaHc6tEG0r
y8p9G3FBaEDfr7Rwk/eIaTpvmjTwEvPt8LS4WmePRiqTXnnTWxPfnBPC7OW6
aeQ8+zPC9Qu8JvcuikDad9NLETVmj/UC6VW6MQZLpYIZwROxjqUaL8dUd5uc
gXm69vWb6JyD+E7a8uNQUNwIzqSYxun2y8h5l6tbGVxKCmL6RmVv3OmLuGgB
C28WgOZHNpe46YDfn73inaF/PGJbtcbeiiT7x2lYVL86rWNkVy2rBAfNwDK7
RAXjJdIaxEo5k+UQssc/+s7hd4qXXMuB3ng/dK7eyV462T8FtZcgbZToX9km
hHsqTEZc0trXdG70Mxo6emwGSjygq0kDAkpgsOkojYEW5VRQX6xI7zigUVeb
uBksAwEP8b0EW6EuINR1H7EGPCG4cGVSm8GlwO+eY9YFlJjL6a0KqUmji+dM
Q43/c2/KNtSwAkdqspa/Igc1BSyTYU1c1LwVLGRx6S2TGJQ2DhfgSFps/yDm
SnYhgAgpOzvvLX/fiPOEbZxJvGO95HPkNyCVczau5MONSJMP32knOrbcNyKk
Ruv6NcczHSFC600WYB15SOSK1ii7oduvBXmxg93DMtWkFw2Qymf+jSEGNIA0
90snjslvSzXIAspegru5KVrNAaHfgDo+gqKD+ZePX2oQaL9RZXKePrW0tZLe
qD+crS06D4PzzSPNRVi5nUUkn/AsFXuC2zMvgg0IMh7LzN/oRo7hTN0KEgck
Zifx4rPbaBRNHtixvnlFrPZQo5a92Hw3OK7G0lf+R4T0sGeaIKYPapn1g/MY
e5aY8I1M82MrCqhHb5JbXZxBKYGL2ZJpK90xcp3UOmSi88sdaA4BLJ4k3RcX
1B6e7k/KFvnzUJt6CgJQ4AxFOa14HnkJFg1/KZaL8kt0sSCuCFmDneBl/WvA
a0jyZLw+1OcD5rbf5TCHTQrf83qdkgyGlt86tLXg25vhg0jw90aHEfdahuq0
LAxdjiYzKw2wziWORRpSSmly2fZkb3Iij6xA9dfRrdWNpM+WWYN95epemUbo
EJOtD0ZFXTEIZOmPRsmcLDczsSgr4iysY2F0MK/VFE3kvgz+C87L72lKFl/E
HzqooSNVEZe24oFYd0PfWWWJY21YqymoKjA7cXPbUu7GHaZ3xXGZhcErxhaa
k8DVcOUB6udoJWE4DtQXJ7b2Z91Pi9DKLXJKdicksU3r6jAApH6VJ9t0pk9/
JK4zYmQhaM7wqGGttkfwlwd7Q2Hxj6a4cYmnQgHNmOSWIYm7RdBd0houfdsD
AJvb9lQGDYv2OwaZ1w0RUO05uL70kby6EjuywwLwTPEzCyT8hdfE8PCtQl8R
YDtAdrHq0bwLATnP9LU6tpkRoogHR8ZOkNDCSh7vJRlehmHBMqhbqa9W49L7
KnYf8It996TBGYCQdSYBfU9pB5lYjUd8njeKTGb76WLfVnW0SLkD1nwEW2IM
NeKjhoFQnHalalnAkZD/NMdGAIiMFh/Ak+IJpENj4IeHx74GRcbkUp1PcxxA
vcHChBb39945xr0xTlQbaZEh7WbPrHXZl2HQkxqXzmYqIkxBPU4WEGuOEJKX
KK61z9nm1hTOObh64lm8n209S/0cZkfYa6GVKtoW2MQnc+uZ1mSzbpUXJETc
MIa7qsVNXrFhU6M4W8rLSE5betZOdaR6pS8e0qqf0GdfhWoyitVpggF/QMC8
F54Yh+Y26XIPGB7/RpkCrD5Zj8+/mbg+jmMJSjQjibwSBnkIwt5jVskgvkih
8qpHpzpjlSWyYDckLKQypRg7oR70rImjBxvsWIK2S/usuZa94PHnMcEYlbJU
7/HP4QYaInSWeB0gvgVMJ5ImgRRRUgKF0iNeo43drc7AxBywAy+/nHXWgLKx
9nUPQTV+irrMF7KGN3YSWzmb/PFJasSHdR5GgEWs3pCmPnPtu6To2VZBAksI
rd4dRuvIwDIlUoDhE209gALOOTjbGYEINNbVn9wRD1b1R1/Jnb5Yc075Eg0T
WM1D1oAZl/tzq84Hzp2zhqECvVdfo5+hmyvFbJGYeW1S4aLoS8wy6+IUPDLM
Otd3Sphgf0FgUi8XjqFnsafSfpt1YsfyEv0kU1xrkhxeTwxRiC+Yt5DoRqPJ
Sk86ojDe0lt9w5ZAkIKJE2XI2eqtjW/Ax5zmEF+5IQcqJD0G7Cs/NvGjOurF
M9h9LT0OCs6zTaR7fBmaoAVVfouHYzMTfrDQbEkikvDz3u9AhV1J2H4mKABO
lVILNxRzvHOf+1tuDFcfw3d2grmIa4h/g96fDYKBtiF1/BdsC2V0NXr51Kix
fNDON+4bmq14bHhbUYcOJ9NV2mx/DRpFLyXBEaiMSuMhoGLQYUv1w9uxjGJj
uTv7xCrexTprWLEq793bhoyuPQjJ1GKXtRcTVJkA9jR+bQyAbfbqkKpXb+O+
ZHcVYkAMSVDQ9xM4BLsweEt10Uao5eZ055vY+ZdTyC065qx+sq/DbPusno+0
4lt2nfwUHVkZZAMWh1lmtpxmX0l7+lRQ1OKshN7PeL6UfuptRSQVeSYwwQMm
6DRS30uaobElBzyC2eRUXlJ1RP83mCFReoZCUs6GMAI2vi6iI+teVQh5mdxE
DQqATyykbAP5bjjKBXbW52PGdydAOzHs7cTCASzIa94AbPoZWhDa9RrR7g4w
aI3Exxi/IvI/jBI0sb3oyGUhEeSIL34i2Tv/JsqJVjDq8khONz/lsEjrUtC6
Ghxh0U34ubdkZ5vIEQ8bAS1xyzIXmqj0JHHlfbfOm6jmcHIEZ+tKnSBfooiT
biJFyyPZ1IKs28eXeJoItIZAAjDgVAWS3WKQGq6SUahf7w0cltcJ8O+5l37v
bJ2mYC4Q5VP5wWJoXPkcicyPjTJkevz3cOG6aU8mgj/6ZGC/tijrUULY5Eea
u9dur7nRjogzB984qcU9UPkvfoswHpaaRjARPl2FQFNDnZTllwGAaCMP1dUK
mRehDibjxo6jt/oZsTHYVfKI0vQGfHF3vWK+0LoAVC4gxpFxSvoC2KQurfPo
nwO+YoGVcJmp95pukKdb/IZgQ3KzIZRBsBu32j2BuhP1alUIQYd6YV6+nFwM
HbNc3XYzZB8HifDqiFuldtUn/GMUqF5UKxh1S5e/uC6gwSa+gR5k5mVtGW1h
oZ9c2EJzMnjDAVdnLo8kIItvA8xiizcVcQq2/rs02B+2aL7m3H93WfjlBWIX
5WOAczlJlisD4zTs4xFflgCpdemBy6EOYjhuHFaFkQiElQoaxh2eNdkF5Ci/
H8uZVE2wcZRbd/XzzcF1/682CLTpORiicRayGQf2hYQnNu+TN1cmPTAs2+bG
PpLnyOU1ZGfR8yL/upyT+x0TwKnOFZUhkkSebzBsIGWMWgRpkp51QG1HSf3Q
oVge1WcYLraUYoeRleFxubHdTQAoFN2nq2I02igAvRET/fZ6bGHOr73ULc5o
WWmaCw2Ai8TW8k7T1FhqBj2fOHgTPv8grY4SGPkLzEb0FzH63fw2gqmDSIRQ
RszLdh+m1FfMMSvh1tA69Xpsg4mNOu0iM/rd4ajyS5+18aY63ejMk/epT6dL
i5/lNhcF2ggLY3NBPhwUth7Qx1Rmkio0xrfx8awfAMnUbg1WhZSzmZB6Pggm
vRGAYkCCYYhIxspIEb4c2h4uj3kmU5ntvCZakqEJRt2IzaRbMhf9rQ66B3gI
vZg1626W6Sx9tFIp7tsNyRqodL46wm+7R71NUyCnpZ94TMrGBx6Qf87yl4Yw
XdDp9biClbLux2w0FIl4LlQTqpZmI0BDnEz0am3lklsH4+avlcrtc3WYUcO+
1SQMxNmusR3zufvloGJMk/DQcHCPwyuANS6MfZxCPK7l4l3n88GRTqcsiSfb
5tSctuw1uMYRlIv5qyGBNAf7hS8BH4nGEoAWvRhqKYt2LPUHiNunTRyF2ejj
eGLWJLnwk402a02frQT5pLXGTbLQhJoRozbAAaK9t3g0GKOKuGS9QqjKLh6U
TbOSLRtznJVH6KmGND80JyDEoifjnwPb0DtcqYGGT+YOW89WtWBuzBwpzDT4
ZiWq9CtSDR6sGuGLCKPw3KasVYjKIe0j27M443HGNtzoh1hTRL+Cy5B7Ryen
eiWUOBZgWs48G/h87uGbADF3bpjtVZSasNexctvp09QX8OJWVzEnd0kApAdk
D7F6dTNzZ4lru1eckKU+gFODCNdrAEHwVA04gL0LMy2B+WjI9vzF4v8mU7u7
cW967iRFdDL8A8AMNXlIaVYG69SIIXoHp3xDtHEKuvAng2twgA7A2qOLKFwn
vhVRiDdEqed7uUhbo7HSklLzajj7XXh53BHWcxKY6A8kOcMxv0lDR7oIBXVS
t8q9YIzhyIhh8WwJGY2+beaaIWq7SsEiJ0U6dK7Y5iZHs+LEk35/EAm+Gd7k
x+QDzF+i2s6gw1tkKteaPR6tkQyLVoWgKdggcgPea9arRV9OSnNvWjcKmiiW
g3vNFZdSzcOozhvjXDtnT5YH8lq4cloMO3GoObBFET5/mP6VoWPUyreTrL7+
CPZrNIKy5FDI9J+OgaRKSZ/cLuIcQ/0FFEOyoH7j3fk+lx99MFhwLr/HJjMe
pjXHV7jYiWUushdLomD5gs2YfSms1HhAJb9Lh5jqaV6ufga/UMMteW2kMNUU
E5t5THc74Hi9Wc5w5AFk8XO8Q7/Ta9SQrNmmlCEHSYZipC+vGh5yxg5gv0EJ
+MbiUuoIQTaeTpvuqcXLqRPhEW2yUubymiVyoALV8UwqPbkg5/w9edSx5708
tLqVNmFwXysML7LpxVMbvBLzf0oLXYeEayN/2H5nRW+rgyBHrZUbGjFqYKJx
fzGJVH3HXnCJuMExkN93H8HzK/ilOs4dYitZqbkGJkuD6QSCfybeXoTsfxkN
zEK71gR1Lk+j5PoIFkbZzrKi6bo4djhB/fLu81RgaxvoRAl4BkVUTne4TbGu
6DffsiwpTHID/fizm9NBu5lWBiZhAG9wS/jUb6hCYLxTeR11wTruiz1a4zfq
xYwaYb5aJ8K+D8o6NffEHQb31O1v893k0LTcKYzUQXV1+aSUUlfOMfX1ZI2e
ONxE7U1nSqFipGV37bJ19onrnUBcbqNsnp7AxkUNtaX4z9rF7C7limWbU+zj
eq4j9Q1Qj/THIyERp/3SseTug9uHW7meNDcsmQrjn7zTwYejguv7LiCtGjup
vF9Rc9Ymkww/wV0YTvmO+3g3zq3rcTEjhdI72z/nP1eLSkbLo8Pj6cUxeU+u
WAgNyQjfh9z6l1kQGL5nUOVdpIARGVgi3O86aiRnT/1wm15UEbdQHkbg/LBh
lQpzedlUmU5gzLl9IhQySPrWgM+9qDCX4IpjKjywA8KGY8oCpqoKkLXcLYd8
YhyUEHiRTZFAQoWWs/SZbdYxvaJIgWc44xZbnwDfwW56KhcVKiro3ymScdUI
Ez9bPGExHgo+fVDpG1B1oAPp7BoNaNSIw8HEXjuxLp+2/ChQGgAN6IwoH7o1
WLKvZ8rLH0pH5YkMMjOO9tVvvdjmhHMUppyvD6Qs6te9BsIrgbrpjUnUHRbz
t2/sfEOiHefzcuMhxl8Q0n1ULJvHmBbpV5L9sEt8YcX765jTWMUsU4QPU+hk
tPh8iotL8L2eiaLit53oK2T5bkm1FLACu96wOrkrKlrpvHoqq5kEWsy3IbrD
XJ3h0PJBUyJo9qoh7/Koiye3bKaEDXsXXRhaQoEz5lcE1mzHzB46qjMnY9ye
BRH+ohmYY7doIi2JhFzSg78ST2s3xry5gimDuSttLxdZG/iClZzlt8ry2Da1
2h7c44rypoudbYEggk8iYjMwgpCPyHc7yNyg1rxg6gSTGaD7/xmclT0kq2Nz
H26w6HM1BEWejjtH27w3I+Sx0wr4Zw/UC6s66QFWAdYW+17/tYq9iSyFReA3
saksOBqw3USR2FLqYaqs/3x1HisbLy+nb6dzzIdEVCBBB2hhcZy+kWhDlAf6
84wYCV+egmcoYtjatZDagkZQ2XATF+mkrN3IiOrc6WGsz4syKrQk805snwl+
TV9BoSdKC9LqghvXF2nIG5WM9hBX0dxivEjX0AqPU4I3ZRkvAAPpr05u9cD2
1SX5//rVy9A3VzZgmo4nwfCHYJSdNYZB6SivsRKjzF6ZBBoDFUiFEGYPVNtF
U5MtiSDnBfbXyOcq7lF1wyWROka23uHxBkOiTqApOsxmv/+cav9ZKrEkQmoT
0vAOg8RJK1VK322UPJboQLbWftfMHtE6SCNOT2tkMb0jUPrQKZMMwB6CZxmj
gtUIBko4Bc2PFX8tLNh25X4sm3c+CClHYTgg3mfvm9HCg8oRc2kfspWkkaAH
Y3Sssap1tOzVtzy/JwVVKMEAeQGY8H3YjSs8EFU5NChTF+MJ+K9NUwO0LpKd
7ZuEIdmilwaXKGITh36cVn81wfx4Fl9BxrFTPslLX9yPopbmGFuItx0UaorT
QDM2bRihwNOSJKIr2N1Lr8bO1M2bnhWj1+1Kg7Ed/YZdotzrFnAv/to/oQjP
FVW4p2c3GR4ANAhHlzh+8m6jGBCYgehS35BiBFavd/qTVHKRcF8y+Tjdzlr/
c8YcbWJHGFeFvRWdf3oklzZE5KvN7LjRPjFY4vXCM3tQrlIBp1Z7sbDpOHON
tGZaZRptXnGiJ+lUTB7718umtWfOVZq2BioiBPcdjbWncm6Pz2OLdv0FNT8A
yWS0lX/FNa9fIBpr+js+qoyYc9Ypzm0EbLdajGaex+KdtmCP7k0StQUIoSBp
1/lyWQzfisONJrXPIi67ZpytJ/kyS4CZssDu6if/mrjfcFawDJtuV34ukZM1
9/mleZpVlFM/cjvXQTfY5Dz1plGRXaVs7Ko992HwuHFpQheiPjplPRUUM79D
MIWW9lo8uPXTkHLaTExt5xMGZFWLTMehJtYdtTh2exR5W/H3UKuW+fqtKjfP
deG1auDPvPMzp9GXXv65qWsc02ngNECCZ0mUj/+gDBTMBG+uKcsYB1XHhEXX
+AF4WBDbsZZiarujQHjpasQdlzQGAe1/jiX3+olu0reFk7Pr3LihlkI5klB5
MDmkL+H9LJEa0N+KakL45TdOdL6NCOXddzNwDp7NU9RFTjHv571DCE4xh3eC
w4IXMa594x+qMGHQgLNTFOVBSWHPQrqC8emGZKxcbadGBQ8cwpbqfVRv5R1H
1kPzkpoW2VFMbmHotpW3HpPf0HZQ/TltCNMTU+qdpAONd2dlH3ioxQABI0SL
Q9kYjJxIjAwGMej46Nod7EXziYcpdmx4J/AW2rrOg7emVTZYgRaendec/D3L
8QKxF/s6ENxCeV2M+rIoYxs/ywP6AcjVw8fZw9yfnc8ApIGpJOpnPMoecAeX
6cMjtgO8D5Nn0PwsLBxffiQOS8Y7f2/dLMYHXoAhCgHU1gFzvpxFXI63H7vA
puHHZLL4/xQoa/lecKBy0f6M2028p/gFQfM6FTZjJz+aypr+PjnZ32XGs3UF
sZj6WHw6+I1eXsPkZ5rVFvYT3jivVOWnVDkb+yhJzmjq3FaFsydfkuCUFo18
TXTNWdRPM70Qq/oDl8ESNxr6OxyHeopB+c4f5Xz/TYiN5HxTd+89bNwSAkNZ
eJqlrP/Na9OgvYCEvAd4pYKOGUXmCb9Pfcr1R6QAEcOGztRNsAMea9Cq+Qg1
HdpMaCuN8gtZqNPHCzeaJ5tUT5KZ7537qwdnFOP26olnAEcweo4cQs2ijfHr
cYqdWw8nO5NCYmNLJekqhLgzSvxUWX+uJs5AZ0EOq556p7+UKvmOS1lEOfTe
BlG9BqqahW8a9uf1IOIwa6OGvKDzyyvzPPzWldMBo+nOZELoZtG2IVO5JhxF
RepzzacV3AHKXN7AHRKHjyV/ItaK3oXATZJSzsUWkFzwEI3+2/SMx91QBO7k
sBxYQdQSuWk+2nX8i8xhNLjVmewnZ09Kxh56o/0pZInEUAkPJeLfWn5H6ZJ6
9MPOB8qnCvWGP6xRV8VKKzwgprTK9RwXWgb8bmiVjXghrwPH6JAxWXWFfZgb
EZaEELLASEM0G9hxldYFFgvQaHATMGwPIydxAWilBbCA7KFvGPOOsWsx6ycy
nW5hYGXosOcv9WbRSpMGuw3nL0yEa6ItavuBjgpmsVpv57Ws8W6I1cNJFxrH
Ht5UY0Rnk5QCIwsw2F1LipOKYLy2MSm8iBMH/abiUTLuOg2neDzjsKyvR3Tg
5eSm+tqWyR4hFZbGcDFlSgxGt1K+nqoTVPoyaYGql5wp7WKPMAkwvHynH2li
qX0RecieAvNREog1iga3bqqfV6jflbC/vZPVH9rsqkx9j6+G1XI2vOBJ0z26
tchnizLTt/PCx551ZnuLia5wZnEIrIVrhYZ3TtUJhZtz0XOZ6dQqJx6VYZdF
4o0Wdc1YMgDpwo7lypiOJQXAFdQI21QP0TTI8acdzCKMgYt5JnCvhmdHXMom
W5ufWPd5a4cMMx+PWwpqKbYRhHav9qHkI8ZkKHgt3n5MJ84daiF2vaBtyhvg
UE77biCsrDV98yPnwU2U5RTZhKE3XZRu/X1cnLH18h54nmBr4zWVD5936r5z
FzC9DgmzsnGxicheiID1m2TjbW9t2fy3mmMEvh354XLBGSVvX1l9//HfAc0U
20ri52AstzPMmqSSa0nkkM2Fce7NNnb1KOJ5RzYsUShbiPtR00xC6GLu3owJ
Cd+tLnp9lnos4D2qchgE5YKgTz+Ns47Z1gNkUUNSgA4RmulCFvV1lG8HcRGC
gjPpL28fWfmncQZNsOGK2W9Rp2HUlP76fdd4EzIsNkn93yBpbKVxrRLs/zEn
mZ6Ucv5JJATfrq9YjR1gCQn4pyz7UpFIWMOtT8X3QmftVu92+S192IVyPf6o
9lKY/bKGZlb5xbLuYuC+OXpO2B8domH6u6DNDes4y7z++IZXHQftkeDZlApp
LXfSZg1YFX89x/gRUL9P44OTz+jmXiMHvl8uV/QDYoGOh+A2Y9i62i0SjUnU
b9uvNUNtPWJ/gu25q2Tu4Q7nYnNsr4sNab5bDvOPXUaIbipZPMMoE3de2WPo
m6XNx6ausfFaUPyT+WQFaFR3bFr6/NXkVoqLH0EWFBw6MsEyaDclfHN9NpxZ
fej/hrq6sENXlCAidIO4t9HZGsZW9s6/kIDG8TGwbwZajvVD4sK+sa6Z/FR3
qP61w67fHEU0Qsg4GQM+epTlKuhJ5yXdaeNVyXo3ZF5uH+fTwQ+HL+rj+XDi
Rk3rC87E+3J0QrIceF3e0LUml4eBA9ICzWa4hU8Guzo5pYzOlKjJa3ABDiYO
yQHITU5VhjlMhj18pJ61sZUH81kmerNEPwQLeVuLN3BYU1bg+DYGIiT8nSeo
mj/KFCc6nN27kJd8ZAVF6BBw1U2CvVjvs/GqSBbjAjzUtmWx5zMPiwwdILeS
N4P1ZjY7vpctgoajZcHk9tGP8bbFyFx2bLsAkAkgohdrn9SkBwyYPHnRloXM
hkK/HfJmbYYuOTmOdfuTiH4NtC9o2KYK6NPek0JjKppZ4aVJD5NZoa4Prrtk
KM/X89218CeDmbwIM9wexa11eMWfRKEMA/s/R91w6SDeI/DHQ9IZdlq9v0GA
5WH7fEJWoMOCiJQdcnbor8JBsYqAwZIbnkDy+ZCfMpIBa6EOJ14ep2qXLUIH
lRn9irD0f6s3W7UROh7swucSl8mDy7AO0LbbthFkE19XNmfyCYs1t2s8LxSr
BrKVjxginR+dhoKdCcPZLqELL3jNkJ26SW9PxH8M4wnJhRfSuNU36B8DZhBe
AEUOry6v737nn3ilWajTsJQxZVdZJ+SJ3yCVlI/2EeiR0K1/pKYgllp+WLFZ
NcyYYpjzQyVCIB5DdaADuwwdRs1x4pr1ageOD4enHfEUBkM4qF1IDbKRQx+C
xfazBtzGAx3bYUQ8R8UL8UPh5AH5zgEgyNQIUqBAXkqIjScSqoJuO8zGrcEx
lwo/wEzag54oc16/LEw0nRFkdrQVPN/RnRExoNjR5dKRHx1lp+p3mPjhx1FH
LAEcGm5BifjT7yIG8VSNFVXAaL39cYCEn5xO7FgHMyez2rP9GBZUWAMvFCgP
pC7rIBQqpfJQUUrpsS4xAhuoaDXLMjfacW+eoZa/sIH9Lb6w5zEJQ/NtD0Ga
PCz9ymc9oJ1ngGEhd22r8cor+x8q/+NlWEdE73MZBMBeTKHpWsXuAE4BBldJ
9yR3/wTzhMx7159Dh9dibX6qS8X3NYCTuPoUUeVhTFwf/uGb6I+gEVh+OZjp
QKgci6puolTh/6PBLL4W+5VJMTLkDOrtzpAgjDpdTZ4d1CReZTbgcj6Q88eH
T87F7ue3C1QEHoY59/QFqw4lGrffSonVZoJO57xBGphlsAznQ9INjyFGajn5
Mg25+TOyyP/1DtBFP/oc8cHFrPImtn4XEK1MGfg/lIJg7NbrZc+phaDv4tsN
AbvxEN7YMK29NVp7BRC4a1tJU0gjXXIAjFXayEba2xJV7rNO/Z5m79zwetDR
AItDj+cJRbkzeOqIdjE/kv4vJ3eNKlE7tVH2CjiT7YNU0Toz8LDZ1i12F2Lg
Ux6YpWkNqJOyP55xYj2lo7rXDDOR1XTOdbwRZ6jntNIeP88NEY7Lu3qvvISY
xAYTSzztQBNyCJ5kPe7/vEIHpHf/mw2w9iWWLzIpdOOT/3CyfdVRuoEOiKXW
Dx36LJYLoOAOq58KLcGCjdoAepAFPxP7pktm46gr6iE2fbTb/OonAVstN+sn
8TtchBWESpQLmfUHQ7xsNgQIDXN6P0W3iCByXjCiBD91qRLc5BqBa6NR4PEQ
/K+7End+JyRGuvXtGJM9Pmf7tC/bPJJur6nbiwpn5YO7wZTLjJhLajTp+CZ0
FeMEmngcgqDXyYViZ2cYqlxnK/4rWhUueTvM+rOWWwXBn95/LlUZ0SW/bSkV
YvkIwI3PVmDJBNjKGGolmse/sxI6Ch7wh8l3q36FxFpBW+HAnlpzsPV6QRNz
Txn87jBYAufIoY0DLy+OmZl+LFPzghC/U0OPr9wMahxpd/at3YDYh5a1WSfU
p2Ko8L6Iy5MA4DrbHoLocTEgqZBs3sgjo+fPwfpSIKASHo6Y5R6XVhmArTWh
dNms5QdefykRP2ZTHYXtAsoInqchQqHSbS1V2YHO9BwVC4EK7svsuKaB2ASm
zlQ/j8RtcgEuYipnQvItGxx2aUH0fAF5SjR2/oOuHB+6HqR3yGgJzSIBW18Y
6ioqvLiYru1JFxQE+90GCcprIReK2HkSONZuD5qQ6AdKMqDpu2SwX1jPxcbV
xbzJcOCCQc95d4Rw15dOvom0P7CN2V6ifL7vy1gQvaJpu085/UbdPTyqBpIN
L/U3JNFezrqvnASqgB9YNSq9aaAS5S09b+11esjFEW8eyzqgKy3xvDNwjfyQ
0MZi9i+6MS1YzgGyaS7ICYfWggCpi1NJufPTqe61NTwQEHWGD6jKznS0hF7k
srX8z5DiWKzQRi3xhmMFUSUGt+b+fkElOKObLPIMmHBi3um+zf/OQUiJzVyp
ysfqLMglVwO+cHgLygl9yH37SzRaNns/0IE2PYjGlFj8FHukl548bZfZ94e8
tGrHzAa7pctAmX+L8CLAd59X59Qi34y6Sn5n1aRMvodVCmylg6mAxw5en8de
bfyK+hkzwdV0CYlWbe8vcUwMYLAwzEeMZnS5YUMQaY7fudkZQ+TtTa4HXrh7
Nvd2Lok0aOg8ayIgedgBEh+UYBfQozEP8+j8O9Haydpd8eygdpL+Gi2ZC3qZ
iH/1up2XEaLwU8rOxHrDJrhIDV9Jz5bnpmwjBnPpqCSDBHbeZUIeCH5kurpP
b8rtQBtbla60CHkDg8QXQebwY+j5IzJHo/G8E8o2dQT+NjIahSpJ9+3gS2ct
DOBt8DPEdqwFk88kgtdyYF9j+I3ocn6nvRUH203RMV1j01sR7tkGALdoETYZ
yJivq8i5FDqlJhIQNW59oH51Xyo/n0YP1nWZwjn+0vfujbrN3pwrBuNXWOX9
URkgT9uZFtxgEXmTlf09ujN4qe/UjaFzHAC8KjVyXJS0fTp00KHQzT0yolFp
zcDB93d4EaNG8p9B+8perQT8NUr6wIx3uAFMN2LmesUUXxSUz74UADazSdmg
x27WwE4KZVEB2CuojN40HfSO4QIACUNo2ux0xudRlK1fAIf32OhhrAreGg3z
7E1zS3Ysl+U3CbKUhdRcjULwsS/yr7cVbSIrk8h8XKdoTnKRiM4U9OpzUGi2
qHcFmKb88RRDeGIaiwYj2gAG3kfZNhD14C/CDwN8GHFNoae/1rGtU2EnX+0O
N5U3tjAH4fVeW5YhnAgltB1MbgexeofvIcf0CEraYlsbnmUSECZVoZrVsZHz
UJsWtygXbCiEX0viD1v3HWhzR2W/7/4Cxpm/yRfb5z7/ZQD9KZc8UL4rpIs8
nKCZDIc6AbYb6GvcupTWWUg/TZ7ay+83FPP/FtPvbRQjAKZsC+0Q247SeOJd
j58YTgGcWEha6wFm6Gd4qAjO5S/TskpMfvv6TeAQ6Lq0NUauGlXi2WJ/gsY5
KmC00GMC/Vfm43CjJG7ErL12vw6fYV7hLzUsfUrappc4Ef+y69gttsJPim11
/OdzsYWipH4P0dEtHkgeTM4T3L6EHOphLn4Ht3m2/GCqSQwjzTbyT6EGJ8Ux
vbuZwvtcYGB4tD+fGng6Uo5bCcx3a5hEP+TEFC1YhKEdVmAapTAgQakQ6K+x
1JMCF2Cud+gZdNiCSvoQmBYfwaEm5CISEcICLIQ6c0gFrWX6J/lNuotYx8Zk
1++Raq+BfYhIdMIKL9aHAfJrHcUM/4NPqIZxwzWZTbtJqu1+36F0pjFKAw6I
AkFgO+yRse23XXJQZGHRYJCIOnFabyiYeQDqOWxoLC3pPex0RH4KXqKS1jHn
eMkhoq5IiAM1jXo9Qs6OerZVMPB5Z/VBfJAz48uTWdxfDuQVvxWpOYv2FbD3
YN73sW8z4AcGiE8qnxG0hBZgeXXyeaH4m9IOZcOF2fzOaqDyg54pEpBCaRni
wbxIzPhJR8JnVRfXdDCQ1UOxA+iZhiiFEFylKQCY/S7iT102/YMjjSZaApGa
foSki8b1Mwvk0v3KuGzmSp+PTX3nJ7U96wrcWz9l8Ah3yXMVeofoAQp5uKEz
vH8FReEctYinK6rTJPz9e0XNQzVI4sYXRTO4O9goTVYF9zlOb4mxyPpsinZM
+f85s8r0amY8T+0K/fZCwybAyRpLcu6hTVzEV8C0yMgQjtH0rSn3YIdsMyGo
CK25cLIKujUO1w6dKSb+aG50WU7ejB6waHDezoM2lmjc3dQ6sWV6+6F0HXv0
GWhnC0u16lL1NFlnwtqqV/9cfeUGQcsl++45lt6LYUCFjMZn2PVs6z5Ai1nE
q6AiNLmhImhPP+Cd5NTZKvAY47tynLpVkw/9YmyO6Achj85JSfx5sf1CqlhI
1+niHUDZmYQgTukEAEIPsi+w2XsCpsGQ1rs+y/9ddd6PrqpxQ/6iGGDUK7Rz
yE6cioafwa0Yp+l112+Ax/LJemQFpTkCj7zCSCHQebhwqEhHLnbdZ9gEfg6v
4s/zgaeuPLvX5yelzpqepHgBRVrPhul+tuGuzpjLBryly989yyOyvLokvkz0
OVifmimljGU6Dp1Mpfgwb5Js3BUBQzIA3qDJmKHAnM2TfgKaBGwEAEeYgR3N
SJJucVHP2YUhzn6R9TUy5yyI60QqnFCTrCoN60n8/ONYx1thvep8jxXuZUmP
yVLtGo69zJ82rsOfo3zQb7DkGKF4q/FwqTPo+IXqea3qc0o2wwqr2Wbud0Lr
z2IptU04mynxVDp76RKnv18GzBJzPlsE2vyyQ4MQpFglR177bONmDtlv3JQM
/Z4ortNZkuSHC16tAWvpDNK17vocwxn7WG9n46PM29+nyVw0J/B3zaTD38st
9ok5Tv7U1/0PEDV1U+IHifxb3EhpKDAkXG1KcDGwibWWQpnJ/PzIuLtJERwv
LY0R/G3+tVbY69Hyd2qQNzrLWQohbUtpaKyDXHzyd35RyL9Hzy2uwMcbQ4J3
qMCaayAlITfamoUbSPu+o8tMgbhubCfF0LvXEOBGuAX6FOusicZTh9mpVhEM
cmEWHNSoUc0S4L2FSkFzCx4z7YQnEnpe8JAuuk5nLdAA0C6rVA/mm14pbib9
1feeQ/lS8+RHC/QYIglJ+uPFkAqz9bnQ7TrvX4R+3AMPbpImBI06/1UplhPy
zqx3l+6wdRWLVgc72GjUU7B+mTTYslW8HXOJvSMg0JoVdiPINp72W4Ekl3OF
3StqDGbGyeCm+84KR3n1pCaFsSv/vQdnR/rW51emrx/9aCWj83Nz3MVesF1S
0F3pjfptW5fL4DRZ9/rwPc5NBaVQX06gUSsI4rjxcWgR01aIfOB8tdkxuOLA
eDgY4+/wloK3diBdaa/6aC3R4hAXoLCw6wEBkXb+GuiEwpEfqVvMx8UzeXX3
HIfCJAAtSwIMPFDzSGMNTOVKGiNZs+oxvVTm7o0fuU7gsUemSY3xLz0o3f1O
w9U74Rv8JXN/N10zOVeltDTa5Voz3VFfYFrCrJMPfpclrcHdUISql4/ikZDc
AqmZC1Qm7wXteHfqO0otFKFa8CJrJftAfwZ4PziTI5JlXvVRoBbaBsv7wn5m
SLIwrXYlSZ348Xbi5EVJCnnJuj4UmUQ6imyO1TPKuY11/BUVB2+85nrmbeQb
nscZto0/1tRrYWSVyKv64Zqf2v/3Z759aQMl9wCdYxw1rIuF+EwvUmoVzYV2
jejqkGeDyjTaobx75SqIwHIVynJP1tcUAdsxmJcjCCgeQxNQNC8xKL2v++a8
LhU/2ELdKJIMAKrPR25AxNZm9T7mWQZIMD4cbxPd9S66zqTGX9KVa+nVlyj4
x+Rw16jm7FmkK7/2by4ezyHV0rivSYoJc+fJ3jDqO24s2/Lsu/8+Yzsbt+tQ
KP9PgxBCl8SK6ySGVG24Xkg2i4Cp3z5Lr3nI4UWqdPc9No3pRxlqaD9LlS2F
MA9pjc53xqaP1NX6p4vWB4scrFpYU2VUR8sezt9JV0RPEVN1KB25vd0zx/UU
d6vxuPoAFb1nrttboSVjQyR1ZNn4WcefkKhz2LYnMzW1+u7rb6hgZQMh0mxs
Famu2TAGF7rXN0lUgRExmLdhbwNcg3IP8WIGFaAUpLBORKCGBjnfszpuz/Ls
T0P5gJoqQRxZp4xgLKW1p3cj9n1XYJqefhhGraC7yQDzn99noH6YQ28hNQTU
7O+3EG/1RFU5lSXMj7WBbZKeVkID0rg55a99npJ/X5ZYniVhyQXUJAizy/G4
o9h0TAd+50aegmBdMbSzc327UU+yHuEslXe3NogqM8K9QRAsyjj8HyD9Ah1g
IZCpfQdFSht8Vat7gH/GApI0+5LzxRjJAf2MRSsI8+Erg/sD4bd4l+5OkQoB
urIa06EMjSfeTIztDz9Sm8Lf8aojLIP0sLYsGQ/V8PE9inPs5mFvKDK9g5Wb
u0jTG4ocULxfA2fu1GyzgQAl8ESKLjZcFrlsyyacWwz9RbzLxMbvTUUXT3kF
FKa+x32AG9iuDI7r4rWUcY4QrDWjVitNfRmUdmThDnnVPICCtUovgaiyYdQr
V2AfttNytBbmrDbDhgHOEPDsmBzXMLc2wKAoBpAewEV+c9YGmLObmK2Py80p
QLRbUQabrkeG5/BdpxkLdVY9Udm+zkZbHmJ+TbKvWW4yBle2JBNygYJv/nWC
D1MuQ79m5uJd4Ue6VKbyUyLUWWrIZRxlD/XqbmYASHTqITQ9iMKT28ITmjqP
kNPG4D6SGMuV/kx5QEgBr11Nt3/tXuSTcxm3Xe5sTdQDkK1dMRRvQgO0GyC9
Zn9KYD1sf2ImnZaSDGFAT9cU9CnSEMgOtjavzbFr+SGKeIWpMVVD8XjLqDxE
12Khjd1E6UoLT8SMhu/SnGxPHNO4SpmgFy61nOg+augy4kq/9KkDNeEjelsZ
t4NwRjxDfmihNChb1BxQn/eRVZXTls1LA+O83BYZZa7CPW3DWRSFeAkHAjxJ
OaI8x7K2bvZo7SpyRgGNQnnO+IeNbFF4gMP5ZOgNYfRkjvBaMuB2OShoQ+nX
qNRbJAp0XMXbwMalqvRxh4fw1y1yf4WJiCOamJkFlPFXA4SsfkIs3W5I/gWK
Ut3VsyuGKFO8SfZYVnaP1xQ0RrD+6zlQJW2obKZRYIcwtd6+fEvduVy/sx8D
k3Pmueqb+jgPhhqxhPRdclaQy/bh8OOtcg65Qd0qNaDTenKacGx623Kr0Pnr
tYbnAMv30AwqcdAnjRJe5bVT+bA4RCXtqP/6M4+myDntj64Gxsmsq1o21bdL
4STi4+oMM9fdIrR9LwyFNjBtoapc+EerBiD3gyvTb1W5g5J9N4R302iNJSId
oL18JMzkGL2vYv/rkai+tYypa6LdSyKB6wyBNXczdyahBj3dEFk5XDcRZmpo
drU9oZFRMZuCWnzzzvccZwWMQUi98WCsKW6kPcEOJaygUls4q+uOs6e2R5F3
Jw+RIVyV+D8YkcrL6klFiaj3xSkMrEJBdwZYQyKn4SVCjYwgc5ADrZ6+KyES
8+T+83Wh9GEUa6XqTGyfEbku7A0EZKrsR31dsKpWPKYn+xoDXEPjJPMBv3Uh
HtHLDbMmxfo8jc6ldluKChwSBi5AP2P7cYrwDqH41/Wm/XBtVzmTXPeJlprt
D6QPjybVdXL9U3dR4bQ8kdDi3AAAK2aWDC2ANMmrfBbzQXKGYNRw7rT7w7tP
Xknf0uh3E3/0uDmC8BFh8/iENmficbBusZEuofSe+IFgh7nu8jfdpKSK1Gkh
f1pP0mdVzWmI/J/puJfdhyUC0OUVBKibs6jNuMhUaQrHsiHZ41yBmJAb/cA6
10OS2q/vO6ccjCXRIxNzSdthjRvWDZJsWEbEe+TsgQr824ahLjtWP1UzZReS
ZoE7zJ5xI58OyLj5ch7OxKRruchjTlSJNx5UKPrRlrXoWZ4qYfdQJkz0/a0O
NeV9r04vJ/ztFlr/nyvez2+ppdmQ4Fm3s+yS2c9xXbpJISYGtktvrSyrg5nD
uQNbOAz4O1ZlUzXNlhZRrxN7KMUUzaGgqkwbcgYzzXHno5pEAscA3/KsBRg8
F6ueVKLhULpD26a7FMh3/QZCzMp0F4GIJIoRwUWVeOQ7Fpa85Hhv/qlM4m2g
f9PzNYX42DIdCsjLnOXvYNekHW6euohgTfHqDXqoOq2AtfF9WJ+G4O/aUm0M
t9sc6UaknnLR4OYGgL4QTcd8RhMTpDzopLF2twVUskg4OgoGucxQwwkx9qxC
F8XyOYMPAWyxbpY3aUE9+Cmf9EQ6GBuLB23wgxQhb52Sf1yV8d39yp2B6DzP
yVErcq0+DJm6kWwh7LhUMHuD7s6I4rZLRulkc7VQhS/Op231aMugOT7qamqi
0jK/bWpkZoLOSvCt2T0tZF1CEkKoy5YMkOgHT1ZYwZJ5WKl7bbzEJoyOw0rV
UdE7fx4MAtO3mrgXrjVOuRz92y1czGvfqDRzY3mQZA67LI0cIHFlAKU/A3QC
quZjvGZj5wfP2HaLEK57pWYgHZMI9zakIh8DDbJR1PKT4UUT+7WVgQarNMas
UrkroF4LR9ssxBH8V7i8Lrz3axRAwnEAZ0+i5GqBeZ3oK9ps52Q758/3xMId
PnHenoHqf/cy4tqDrMLmneeT5adPzfinvjlGy2PUYE9QdnwGA078RSKG6DbE
qmVtfTlXDfpD5I02AU3Fi7Farf8dggqzSsdnmnZHnjbjycWoea3p3ZMMdMuL
W/q3J9/kYAll/CWG1RzrWFy8OWWJzaq2CwQOoOzXUJG8SOAKNfSABNamZYUU
tVhTWJIh7L2JC+N0vG3VnY1jax6rrwlV34ePRK9XA46fwPoIGxFRdlMJKhbP
xlSiCroaKwCtcHtn5kdAYCV/qFjvbYt2eB8+6rXqhEqX9MXoh+eev1814hFR
CizNIlojD/Z3ZRZA0cYn06NZaDf5x19Ejbf3wTW/yzNG3p6qx7oL19/mXnjf
8Ls51v5HonqCrk5l8jyGz25Hu1+PXLTkhgMwo7jsF4o9rkdMDqATtglIj3UK
El9NDplc0c6zUeaMbOwrKOkfVqdzXhBYzYx0tnIRvMfCigf7MIr32XUPCJht
zghseKaOwqmruBG1BQUhyRmDfXcs8F0HBMCwGUhXirguuH+oQyM0ytR+PiF9
J2IYfGLjYvMGouYJEx4ucw4yAzYOaz3rJtNsIQ7+CcFAvl1yAkU4viwfr5PE
oriSxrR/ZQprZ5HEPFJK6zKh89FE9+J89Gtu4l0Ic7wcxji5PNMwy2l0W712
T4ZoiO1ZlR66XnogRITQR+rxiECQaxhwCokOD5f5mVqPDVZbHIX2yH8+uJHS
25MapKYtwWoK/9wOS1Bc6toFTg/KzFOCN9Rp20i6wV3mcCpMkpAkJoWiTgMQ
2fA+HTP1npxsl0P3mMcmBAV9CPd8CbDbe8uIKEsLmDMl0aIdaOFRma7cnWnB
YkjrSab7ZcthdTy6euWuSz31ldPMNJPnTRosSHtiWEch4AGhGgnH7EfPaDRb
H4M1XlPW9FYWZBs8aJOC/IGfw5yqZfckucEPMZdntWuctOsLDIKHhccBvm1n
Pjm84rcm3Baud9hkgFPRMeLPeGlohezfLzUP+TkwgXqoSN8JJe/+bSZxUtIK
idhWIkk+CZLPP67ImPSmC8RfG28ZtU4CMkNMiaLLcYKtgDnLD0my4v9dWzw8
Jjq9TVlVZ4R5oawSXY8r5hHy2bQVraGnofEPlQVi5ovHMqCRIN4a3YBaIdYN
/VYaSSSSXtACPfELnNEFTuhDzcRITZ/FgrDT/XjzEE2hutRRaZffJTPFKY7G
+tDxJNXnQkMlaHXRVLbNuWkKuLwLUwYBbA5w5uAk204Uko7wtHSyWv9UDk2Q
/Ut6F3TmRvPNoe6O/uzs9sZO/ZgpmnC4vuIlCtAiN61mTpRppd5QGDMJS+n2
HZesUwVnUIPoW+IrgcYIpKqVH6GpSWpuQw9kpxljqlD56Q3oF9x2pnIjkW3a
GaR3/qMwI78iyLdFNlt/v7DSvAna1TVEnwkJP8c8cz031xhdHN2lU4hEoAOz
I8TjXjZy1TiLvvMjU9bQO9t4vxTRP3fv2Y/47k2nc92eUgVwlBdtAfPQRIaD
IuVxaH+I3Sem39LMqBM7s7efXSBlVScDe62UvqMP0hUef1piVSa/10wKf0NR
hs5k8eK4TRQTABmqatodRwp6iKYuptSOboshWrVGqrAOPwI/KAjE5QMfThLX
XI7GQHfYgnWv7DbCoSNLTCH58vLwJh5p31GLhEv9t0AEs7OlTzVD2iDG0Kza
LG18lwtJ29x9CZNCOy13LqUinaCNCJu7+X1sLeaUsOCaA4GUOK9IJLHe3OxL
M8vjmEfxQiC3LNjWJT6z+ecunqFLkELVQFo52JFyglwVmchaCy8BAN+L6DDk
cTGciFXPmyHLt/yLN+gcWLVe1bTpWfof4XZy6mc2Q/bquE6rqnAMo1J7irDe
UagLar3sYGrJ0FuPJXZWCePFHDCZ1dTD5ocjgmsMVsBvMcKcPL0bMjjHWvQd
B9g6UB3wWB5yZIiS9KbRNsF04DgrF1m15xQUzxxmqnI/6FGHmMNkV0FuQ81l
7tuIScrJ15EFTeORcBlSvcCooP9Kwm6SK5Z+82+zYhluDqwyWBqlxdopSPcb
yaO05U+scF7CnYkdbcclBaYI70iDJdB9f8nW4AYJJ3QqYrTFwsFXI9CrpPMu
ysmM6KmKQunM4VoJZFluJZX3R2zLdPiaApirMRB5uTu+cxd+Q1twePzuj+h3
B1E2QuA7PylRk6E8iWOiLf+1h4SsT1Sv7XKpZg3iU3YAriz1F/ifv7raLWhI
y/oU1Bpjej44agL7oFCkNytx9UaUZJ1Mnew0xAmpumdUXKEAAVu14c4AtDdf
Mwfd2EhFReW43g39CRs3nlfC1nQMNGTEuetgxFGVLXutzsz3B78qNBmq5vbt
uinY1asHhm4tC5K565H/MkRFrqHqYwBwSmcbwhI9z3d53959gluSZr4YhA6L
DCq1y8oxq4FdJQCUfaN6g4/g2X85cm9ew7IopNFawpg3GkulFWXcKtPgwSbm
Ps5Txr3O6IuoUFJ8Hd+TqD30Ks0kkgtHJ/97Uw+XXAwAmTAfdy6A0+5UZxxJ
ACTG8m6ZgnZ4lTfchlTkuF7U7Uvm00J08PrMJrU6UCOl1uJ6XKaEwGqpkGaN
QWZfWsVL75r41QDF+Nok57K1RiBbp/Fq6KI/gD6NI8R2gpuzMUrIlHaIp2Uh
DTzL6HreGSX/cnM5Y77iQfk6/R3ejdBBDFElenpQJ5/391/Nue2uuQXQupXk
FeMLVV/6Fvw3NepgX7+RXmOCiTPmx9ccwTHLWLCUews3Xx0n8aZFXVpSMWdu
Nmi+rUSBocenXlhPisCTsD51Ff7oTP4C1EEUvDOi4+FCAU3CAGo28UGYEFVp
me8tFzLd83lhWwI6Zh/vfoTOiGS3sRj+SNgtvrfkpADtEsgvfIE3W9b5PXtB
RkjtKAp1X8Sez59hsmMOO/t+HZq+eVzftRQr7ajLHmUNhTyvtQciJAOiC075
mbo1beEDV97F9MAt8ZD98q7e2r4aARwtlK9dTOZRQUnzPgH29KvDq8WmDEzc
efggY/NYbON2+nvthXeHkNW9RvEFO7RO/9CrMJDEdXaNjbgoxi+2a8iOLOgK
EiMmg6BBHn68gBG6W//EyGDY2UkUY2YZ22UboP0WtsRHnaIZU97Z7CHPUMmD
3asyt1QW1qOtSOpeHquspxIPkTyh0kPWvWN1Nck2uLC/fQynZrpm8D2Ti4YR
2ClLwMVksioWIEkoCOm0UC7lrNdW/Jm6b7XH8GacTfaEbo96zx1spi0DZqqR
yrGDMZT6u7WR0RMsnRKcTEj9jeY+FfAm+ZsRPkYMIMiL7l2wuyTbnlT4/jMK
K6KlyCBBma13GPqPOyfd5qIoc8Uw6osxkM5uFKaBdSgi26diNJvv8ZJ/69eV
maz1uCOQWadgUZ+zYceqBFckWHqPcr4dZpwsUd5BRufNOa1cq5vcklwT1kO7
vdPjRoAHUhGSRMaNy+sR7s9Vlzp4jOeBaydSlPyCeev9H1rMGtrUByGFukOX
vaJk/jxTOZvu4Qb/7/BEBChc+9KAyBxRiFoJETIn/iOZy2IRHZuVSUoMAGgo
Ki4jAdN6pEiwa/BAkD8GcL0z5IQ962Wuay/KepCmyqPy1gayOEUYMhM+HCOH
cXfs7XBCbDrqqI8mqZkq0CNSDIf8ZcXS0Lh9U0gEvuYKEEDt6/ba5S7jnsrO
IEkidI6mknsOD/gF1zg1LAnNNY6ztwcskMm3+pPzONz+fTYUe/9ejlEzhOw7
VNZIeeHpLnI/pw/nOQYHCQDiKHZXUrhjJd9LUiFCQxE44dA/6eq8pUMkPbVK
ewSDcIznrEbzzRnZyH4hTjYLR2OOWaGH+ftlzkH2C1770e3WC2ZNYI9+NwUC
B9RLglQUlOxSyPHrUnZtog6UoeGpMKndVgH8m6WnpTth8XWGdQN9Wixl7T8z
eMZUwYhOL0hBhSWHlJKrzt8a1ahTGF0O2iZJpFwVA+OlyJYlAcISzFaOCMC5
vSOB7i/JaMttDxNrAx8SlO4sag5jWAKROQMaGrLoB+Gk0uPCBPgAXcx0DzcW
13ryH4FYV4RPKMbRPuaNzTWfiHgshoHw2pjfiZfInW0bfYoQSLfb4i0nAh1b
VP+BkkK74WXzGm7ZU9fjyj/q7VwBmCw1DRV6qRdWp8Vs4M7jll3KExGsE9Vj
QomaxVLRpNsqhyg8Dp7578YaUkE5raW+W0JQZTowAD5aioeyBiJr9F7QDt0/
3ZFIymrc2NrqkDeLStzZZuc98XODnFXfrKPovuXf1bL24J+s7ilN4jnAQt0k
yi2RYqQqUotjpIWuLEEL+iUVSaWwh7NON3pCPAapN6yKt8kJKgxjLbTXLMC8
VI6d7okukQUgDvIjTSGX5/V/SBF8ZMT5Sj35i0HYe94iTmtqsOWlbkB8fLFg
AQxNrxPJ9daP3JKQLssE5d18g/QFg/WmaKo6hF50lE7NB/51jk6aMrRRCjR8
efYnIajkUdB0B6NnVv11a/FAEmgthjf9CDO0s67DjaQJslZ9eTCiBTmJmHYQ
85Cq4gB0oXBIz+LllfNoQq1PgXBVF9RAdkGf8KBLi5bTlkxjNb7ovcmmKhrF
Z4OvggwUtWUUT2asSFhX7ld50Gc6o2re4PqkTqjBMfQcDzH4t7Y4U56hxCWN
ZI1UAo7GumHRJrR4bd/4eV6PbHaFI5fgj4FD5PEMhXHXoCe82IKp2DWfwe/w
liIyguLuKLCvdps91CcDto65wogh6yGN6qk94by593bdQM+e9ifOAICG0Hrr
H+uchtS1n6sogDILfFJ8clm/Em8lg/QdkLRenu0cGFxaWbVcsVhka4ue3o5t
KG2+5hmGvQKJIzmlnlR9fFW9G+Vs7c5RBhfb1zjXo6UvzP2UYdACv74my2ic
1CdlvuCcJwohge3lnTgZ+KEID2Wcr8wKz86O/paH6UxMtNCcPJTRk1G9XThg
Q1xitRNgAu4Yj47LZo51iNZZUWOva8AlQhT8/rpkWh9yj4usNJocv6Z9XDNP
TuXc+zCG+rP8tGVnh1hmUdu3LwSL8ZZv2232fFRWL8QuHKWqXWScoGY+OQ7Y
PnlwCLtGB98kK5IYcOcAyTnQc1Potd78ubm7zLQ/j4RtnZlGslIQBILnhjly
3H8rZTF+3cptSHUTTWxZvY3GNoxzt7fP6GDQBHPlRT9wOLvuZrXEhConNH8O
6hUA6gzyM8gUsxvpfbux5CDKjHWJfGCVWdcWRb6g5L8MQpviIpnL6A7F4q+x
vjPQXqWV5fB42/EwrYOvhSGQq0+gngR3Wk04JddFBZUzqxIxt4gUM2de6vBM
WwDo+LjtGi1Z2v57I6fidumZRSxE02TaSl4KLPNxE7751lSPi27CDxxgGvou
xoiwDSIcDQ7Hs1+OXq4RdfgZnfMekIyEn78NgO+mHB3yQx4Ajjv7UCNX+l58
z+3HoGfDzwwJp88QNDw/+DmZpeILWhS+wGo6sNuEQ+oOVJNexTTUvF+T1YwK
nZJ9/3WemeWTeW+Ybgp7amg4hyo+okzcJv7X/HUEny68chDkO256g5ZAcBrk
6Gs/7+hmrpXjbu2CLZ8xnTBgeQGh23hMJQDtNoIRpxhnFm9rRjaw/DHGAXu8
S1YktXDGC5pSDuW1h81zWZOPsQ/AkT4iS/LJeqWBhlvDsyufqKuu0zWk/j94
LEPZb4o2zTE2WDUWFyCCxjgqfkHAHdn+7RgO0p8yfeHl8ah1sNU7zuTyEGCL
4Qi9T/vrFQ+WJV4NoBxviS3TTH386BgVTVJ19wTuL0odxtHtS9FOouDTPoyk
ONGxxLvMTau9lFG57jI+vnLKWLWc747SmhUubzydXg8Ezf9MRLCX9bZXyA3m
KMocqQTCNANtrh8uN9IQF+PxsilnpaFCMM7mqYmYwvcdvi8XW5Uz5yGSMCT6
H2kw+y6BQZ/7fGL4Jkxq1+F3xv2FaQfCFo5FWHkjaElfs+yQ0xj+tpE5Jbid
z/J+IBoNkzrIkRKxLWq+tlkj9xU1HPt4ifRxr2AXzfK6YZTYNAM+Ru2Q/m2a
rJNLwIQpfeqQtiP6Y2hl47I7r/ucFBjI9jioLseMJeXfdnW1KL28kEgEB8FE
1NrJassw+h54GT9YsEszmIM2lCzYWc2MdKWyJVvQ9jbmQ5mCZztAf4HyP/bN
MDf6LqaDGmzT9aYVNoOPDHYu/aBoxBrHmX8Dm3whULO5staaBEn506QrrSFT
mI8wfgiySItim3t8Xujb5cp1GRDu1Su0wvv3jwllhycPcq3yBP9EjJzgeI+m
qC8V6dMt1ayZnR/coF9Sobyv6q0qZvxFT26qKkAkdQA6CUOgXJB6tOa+RubI
4j6T+8XEROVcKbHITPK+bPyD6c+Hw3X52beNmAvaWimAbt/UZi4gt2lJP0Vq
3AX9aA7emqhxjLcQ9TkOvTTe+0fMpbpftS75XXDBT0Wcus3J8zcrxtIHNmkR
5KblCLrNWOsDIDlIH2OIX79jQdgdSPDig7Cad9jKDZzEBZiSVUvZwIEv/cvj
DrFjJvAsC9hWsXYxKDUaThbTzI7dpRCladqpTXEl5ZcoCrHfQFnaezCHuoLe
WEGnYwxsJbsRtqFfzM9IS92y240PLCzUbR+ZCUA3JHYfL1lgXkD4JXrsVLl1
D7GbCSI8Yzi/p1G6SVDRayxiXcvfT74IbTVKJVg/DhhHhjbPnxXU62lO+VTD
CwCjXccLu0GHIxWAFpTaBCfv8sfV1JvITzxEGIrgo7w0qClD1B6QCc4FDl+N
TYJgfYNPoCg7LoC+9jhUpE6NHcizlZ+q1QHcTcaDJmBdYvMO3oeFKMZt0VwK
SFI3+LM8Si1xN3M6svger1Uu2n216k4VOnwtF0h8CiHVBMaKtX9+e1t9ExOC
r8O4IxfhRiJBm/+oDy3Dk/nWCzvJC+9PGF6OWBYKsi30zKzCg8HJuw72UjYr
sjmw0xkz8HdNx1wp6vedxS4egRTJcgnMxsrYbPwrs6ivq66F1I5el0G/oZjQ
3UDj79/qKCVu/xig06GC/k55jjDyARL/PrPxd7WgaSvBpiYYFJgM4pkhzWUP
fLG9j+z17d2cb4KwAmod0hChJdaSYeF3+ZUYqYulR5xdL+UcJtc7hM7rWpEL
wWxo1mM9inudpNbeRjVAtc9BhT5PviB+RatVrEDosnjjDeSp/qqGzR3Xvisk
US6hNZR7Bp+uY3Ir9z90hRmpfdEiTEdWS0+bnlHCva1G9Bqwi2KOe5+9C/IZ
DpfabV8bn8C/nH3y2fHZxdnmzGjLbV5flwG0Pu0jSItm16eiPna6dx3fHVsq
zUPtu0GWNqxg90cN3vk16I3TgCxGci9NP77A4/ngWgUQq22Pxa4Msv4EERPG
AKBkQR+hNGRX8s9/Vc0yH1Cfa/VcMCv4GlCrwhiF56yL1f8JI4NJr+NrDXaA
zEfxGhBG3Z1hcx1oPm8FbsElAp2syaEeX6rKyQD9B+21kLdtEUbA5hsi5m6/
tUw4PZXwIpi8oIjYHucouYZjjA6jSuAaJ2L+kjZCwC3chqHe+tLINJQzKIJc
xn6kt6PKKWmTnUDY2AAUDf20MlGokbmE7eMQ66J6uLQlPqg5UyUEt+StkZer
pULQDKh5AmxjiucO0sxnKx8eNEwgSrVTNKoVgxWe1rJ24rU8FIrrH+u77U9h
eR7Ou8Ri4ZOQiEem2nSNJTlEuiVf2f4zPOXAFapvASnmnzCSEwFYlc47OigR
8hioWUxuaVONHPk3pKeUUSA39Wuxfl59YflL1MDd0HkOUjdHs4KB+S91ytwN
LPNiCt/UcXPZkrGPO0UQSRGw2KQf/X0e75bfMQv8w6KR99aAp0/+5zciDanK
WmCOpxX4yllSTOUKyPf4t56Swu/XGZeDW6QmZST9aW37qwvUeoRRiWOTME2I
6KL8vIrZHwsuFP76/Q/CoTTpCPF3fEXf2/aPNc2+CPordMxD788oFpLasSY/
pecgciLFe+FkheiaKPdMLZxarnmOupkcNfK4n+Lw9EnPWGPW950byrhC4aPO
NCrwoQm73JKh7jWGiznm3l0n8U59lKLxGQmzfeAEMruNtBWS4m0NqfvvIvxX
AHMzAQWDRveudwmAzkZzS1LPigCO3xi4GOuaH/Vwzhc9GgUziAiTuWezRT1v
cP117tPd8i92D/ZJLopvyiY7s8YkyP2Ye2olR0VdCouOmjoBYU7xhTbQrzbx
MMWbuLPzinGYQHMdka0qX5A5qERUlsNJdjaFtQfSxMfwckJlkgD6ajEi55T3
xbd2q8LTmn2a1OkMRNzda5wpNyyqV5B9ScCxsWxOC1qN1xQFqJlmN8PznoGA
Uu3OoCz+Dh6mx2o8ZV1ZqTJAf3IJbc0BZlFje+w9cV528EOtAOunRRkzVLcJ
Zq+Sss94SihdH5KNXXghBpv5YGEcVkDkKl7Fr7tS3EsgiA10CBh5W3awAMNk
mAHh2JzP6kyCp+01ppKcTFA480tfeO7E73mM3MyH4fbctTvQtHRwesWH5mzA
ety+JDwJDfeZ6T4T90mWSqu3OfLqp2hlDKdo7yz/mJZKvv7jrce+lBaEyLkg
0V+t2PgBxFNgZf7m707LcOu8KmaB8SBxbI2ZbbMgVK5r31EUpvGgBwsDL1rn
56fUI8UXtohZbPZ+mrm9eVqNPZYYC65YKyCuLwcHVCbclbdE4ZPG3YwXt3mG
wQyFczhBe9hnxdjVkYqg0gHjbISQD4gCV6lVr9THHXtv+kWZoIlhzt7aZH/b
1ok4V+1+1gcH9eEuO+Hlsn/ZCBqLInEW1yDio4YxE71lIlwh9y05mfrLl2OE
NILT+5RCurFNFwkCt+b0cPJ9B3lvUZNN0oHDNhqweXZAP8qWsHqBkGIWPBgX
pqJzw8urrCA4XafAsVI37pYBUqZ9EIO0v/Ac4vnj1XZCopN9Nt3ZaoiXe55W
EfEQxKwH1FVamTjoPPiTRibXz55Y3Gu69w8R0TMcXYmcdovWcxJ7d07pltPs
dvq/fK/K+/gapVX/KWuXlJynmC8uMqo7cSxLADKfJTxTJjTD9RwCXYtyWZaF
Tn24CF49++jay5Wlx0jfPgQn6PFLPqmWONT1dFc8gQi2ZCGhK2wIsyI4G3ii
+ClUgS4U16e1xC8GMoZrY9WNbG3omg2JLYwEX6KAarA8FeUAnvF5OgHlU9jG
ckbHZoZPT43NqHNvKAa9HqVP475xgaHsjp7EjlyCONdu3756D6YNyA8idG9v
4OvTQY8z/hixML1riQYXNBs7r5lsd/bkL4Ihy11lJfLjjXtVw/TeWlFnE4qP
UFKHcyX9z8L+IFjnfiL0AV/YL09tbOr0aAQVQ6SQafr/vwREnsb6E1Ud7fsz
us7RIh5+ahSGHPAR+IlkZTF/+R1HHdWBFZ8CR5DtmLED/YeVZemF2KCwB5SM
VIKX9+Nqs2vgrZ++z0gRKekzJn1vw80Hcan2YD5KKTKv8n2g3XQsLXO7G/sQ
hZlDUlkBZDYCxH5vNR3A6JMYdCGYVNqggHyLLEzaIV0EQP0Bi4KUiFIAj32t
QDAiS4yV8DFPSmB9cRoP2itZ8cb+5cG7Bh6NCcWQy8hYgVjQlofbKp3sGpt8
SpsLlb6l1OYwebZHKQx2IjBwJ6VTNOpcYA5vqqSuj6lZkhS+NzbDzG51Z1Wi
mZwsW1Ku15c/TQ57QIp4X47/XO4+ivpJAmOM5/ig1qxa//L0K2ae6b9CyRCJ
fPtSR9Z7cUE2aGcRvQRC2OaAfdXf8p7V2+INUkIaOQ9o+ThZbW20z5v5DLPt
e5WZk0c2OzpqSrJPFXpm4QmeYhS1kkxiwbFjhWXZcixlXRsutXADEd6ZAWQB
XeevzwcbyLcBNAkaNXb0frd7NC9lkjuGdaFJUp8M66GVahOwkY3Ii8eIS5SI
ZXiRmwms1bd8T9Zi2xUucdADlAJvgLBBkc2wobiUURJmTj2NUno1E3rI0uqb
a1Qif/0OMlqbIE9DiB2E7HJf/t+djXZP725uh3JJ7GSVH3gMqXpWx3K/h4IF
+VznCgICt7jq2FiKoAOFjpXefe24JuVnkizPKRoYfpqihp758p483VwmQz0X
Xna9Ggn8CRNPn4HsT+hB4laQiyhHf88NpR2TrSc4y19okl0z30C4zeZNpZGn
EGmVVaVgH9IX9NcXVsGixZxxNkliDdAvoB3jcxO7TadIM+JyagSUDHbuuXbZ
IiqCU/HJDfyRchmK0J3tA3nWTD4h6hZvISBlTGv1YPbXUEQpCoWVWpB4Y8+i
GjJppf2D+S0Wg3ZaOec1XxOnPGVG0YSbiiy9cfcBQaYHbulzvtgjWejP2N0l
2a67yziy8tbD0h7Kwugd9MgvB4ByL/uXuV8i9+q8pJZ4DiQjozC8T/VvnL03
cjBzil9lNh/NQlZ1jQaWDBWSsIh9TxRKiwHZyURmNJY+hQMf6Dv5rTxi5A7i
ZtYw0i9QDmRQofXlqI57iuog7UmrEFitwMkZFReFGmipBddQi0Rl6YktcUVs
jwfJo0tXVtkLkDKPo6zOGvresJigHT5eAiui1kMqsg5l02fk3LNTxjvD5N+N
+/TY/jxjz9VVIJHjEaol2iUYEaGFLq+B+CmWnMJHFt5osDcvR4IpVYjKGfe7
k/F7j3+QzArSb5hpdRlMEajh3t0qK9rN2BrXrdCbkU6A5Sf8SU9dPr75wjcs
/vmjl7+1NVAiA9UWdQXa5RRIaD8KXRZIteAeigi68l1qn05jLEQ+7T0kzL6X
k9Bu21ixSCRGw2Qo3RWs2EqG27zo3luB9leVUIQ420E+KNFj6bXoZwha9WiD
Wod7tlYWUa4BSZvBZax6jVi9w/slXUvCUuY06FUctke//ZsHsuUQDdxNhaop
82VY1Dx0MhQEfgU2RGRQ5bNcnqqQ4BSU4b0+7ywDgvG9jdniqierwlO9ekgB
Hjp55okKcuRDVPcR1hCaO/7cUBJY7b6MMkbQoL2nAMsoW1IcbIZvZfht+QM6
vUB3TTKFNoBUPmp4pV0RNjOpFmqHdWIzdQ7Kw1pZUo70vSz5HGl3ZC0ihrTn
CEAz/c3mirFVlsw4rDn3e0fZ9Se4iiJ7a6onEB23bd/PI03lBU8PNrog3d2e
eQYivrYqsKKt8vbmbbDm+v9CXMXJgeJuNiZXXo3Zhx/mj4ULbimZrjBAtWzm
DK3Dg+OP6d5h0lifII3LIZUnpPU5TLYHJqQ4QJe08ZuLIgrZxjLQPXpS55Qy
6XmYcjePne/5WzDpkd8N9AAoX9Qgznb/c5ywX8yhOn0tbHlPe9fNAQuemfoQ
dxXN+LN4TXJ1Y+VX8/PimmkmjP1qpExwT84ZvSEB3jlqi90ORBJw/FRuIZ3u
yNrMAwvWE+99GLkKQaCX/+jNujx84FRiVZ9j4T8c5GilaAAaS2SoNJ1+AsYB
V89iBlgQ0r69SVf9daTQMsGcBiF52hIyfEZcprVOvNKGT8fkpKVLIto7ebw3
c3KjO/vZdpQcTgMG/Spqm0G40Ec23tf6CRW2m7br+fHcvmYQeX/BmJo7m5fY
j38Vn6lVLZpQDWOSno5gHH6KcRAfwYfRqgfjIgDZrazlJwSWDf3fsIrAOPHS
kUgmNx59jAVFF4fwTJzhkNV0IpXbJTW+BHsI4bswpoHiA72aFeVHac/1ivVs
4Kfz47YlLVHW7GckgNKQsuMFCcYDmFujmaC5C3C0k1ZGNVqEomTVYmI/Ekr8
KiFk4Ol3YGG0IBxSp6Y8PcUNWfd1jf9fbJnljbD1P7rDoIN7spRpdvtwdtS5
khVzqpw6AVIGhKBKUwRBAPmTq24//YNkMgJTUW1bgrmIYhLY25G53F+URKd6
a0MBFqX19KplQ1po0URxlO31G2D+SrRcdOPwpgMBMPdQdN+4QOcOJeuu2SAz
/QBDRM9PApy23GbHhPUJf58ssGZejYBIOQ0Y19G08u/Q1YCRIs55GvAttzKO
Ed+O68ocT2Hb5eA6W+2sAlfzOKZk13LgymAtTfPB94ZxCS9TPEkan4fFAdFF
Fi3pew31Q0HYpZR5xRGnR47weQ8mjxj2ZmU6VNag8GPW0WUArx38vLa1TlVa
ov6qvymvGeLocVyGeysgXDfAHPYVf+TmNcGszqhPAh+0Sq7s1qd9GDxCwY/k
fYjNbTmn2a+E1n2XGG7pMUVjhNPUkCXYVCAmZk4qNqbfn+BAJn8s8a5Banrb
dyJteOQ7+8FCrZ4zhpq7QEIB8w9ie93Zd5mRRSk0Dyf1hw9Y2bNZUKca9KpF
NYznVsNLsQl79Dt70uhzE3DDMwpQz7qPNzghCN1Akr9q9tOLImM9FqGOe1vc
k6+SshEd/MMBHIBXLK5de8AeBt0x8cprzPag1MclKWW1pK+gKAcrXt+eKtK3
WwqNCYnuSwncqqWlnPTcafnS9vripANlWi6jiRy5hK6Yzp0qr8+ZmaQkoMrA
YZR7Lota7mx04S6boCIdmgMoJzFUsIJBL8KSpuIAcKQ3kjpgH/t4oYyQ5dTK
sklSFFTKlBUPJI+QneQEkYGz7x+Ub5o8pmsuCMYVZjhmun7SIV0VkHCcvHno
ckwRrMZ4kbJEG2cKEu1pVTV8JrRjs10ET2ZJMbafCLEHgGqYASwZjVBB7rn/
2t8hV2FP8DFJseJWNjFYWtG1ISo7AwS3C3xHdBRyZFNxCpcQgcrEkA49CS8i
ygKvbQ96QoKveXqD69tqly8zF2w31wu0R2k7YHBgOT0n42TzZTDqwne8SKFi
wF+NXP75eo0y9D8QhZFmgPde3bSKSv92PSsKQdLdjfnMqrEo2lDNVUT07+nI
PopLnqFb2kpgbIvrxuGjXnAnbY0KAgF6zy17rTGj6vN60Q7udw6oGJoi4LjA
epH5rGwqNW86JHcYAzD8nSgfuK5mRL7gUAMsOzK8+CQyxc+SZSxuU/b6US4v
SEUvO/rv8RyE/xFKLFc3l87Yx2W2wUC3qRHZifHZA/W/Wh8en4lcMUbd5e2L
sUP2d/JvY1bix6/Snc7jjaHDp8DqQYVrNiqkcz628gHgzg8siAy5ErE1j8S1
q9UuEy+cYNKNc8OONf3xalWGp5HTCfzcph02xSUbJy9Ao+cpdQPTjH4rJn0S
W6T0YcQLKh1PHIuJGIHD3//e15SQEhrnVQdGKInUv/Q0DIK8wQRTbjHB0djR
ISVrS5tprgXIVrp1QkTipZ5m/mzEJgihh0+M6F4UmVl2YvFQh8O4L9JM33tg
XfmL9IWGaf7CT+qU9K2qafe+Pf9WHLXvCnwVUTwh0fC81fnVGFV5YjvZbSK2
XcTvFdK9xqvEurmYgfirKCDMCs1Acwvl4jh1ibRUd99P1RnyGpLplN542ZiO
NQA5hJ/085D9pC+Xs5BkEQHgvRSba984B0qevmKnmQf+cYp4LSvB1bj71Cb/
kjbt2QDii+ZaSX3buTzovqXR8PylMiALGe5GkEBWE6SPdkZweUncd6yA7Wet
/9MC5sJEX7/EhQo+aIDRGeP08wUKJEmJKNc28k1ptlO9br8gc233vqXh2OOA
dhe6i2JNurhYNKzx8PuIJR3qgMXKNpYcB0ZhHx8MGC8rlPQnNmFQI5p6ORg/
4eC7HgcWTOg3WOJ1zlD9iLXSaJhgCfxUkOra9yWzUels77M8O0LOCRCYurIj
yQifBd8ygJT1B1mICEQCcQlFDPzSTVgtXsSDdBQEhhlor4oo+FYzunyXxH9X
p7+PxbvT4PCYH5GaznTkqaQI7qz+VYubNG5vW/PoS8JsMvXQ30UdgbIQfuv2
sffOSiF98QEzmOh0tNrsz04JUzKMQFyMdK1jO+OVkt8txvxBt5blI/vs5pqv
q/RCPveq9QMLsUiexVhD32aiiQDdUgjH5l64gP4cGxhhpNDCib897/wUqDKb
o1ozljB5MTU10JSuKUmvInUeel8z/rsXm5bvliB70F8F3hLkBB1st8IjrHBr
96ulKx0+K1gb2nKB5xSgAJ6nj91KqTI4xUwvNs1fL4Efvt6K6Ci6Gv+iar11
WI6QnO6IRU0dqXtE0r+LJV6pbxdu3sFZ7bwdonug1SUay4HAFDFROICXHuTj
1bzaxRWNsZp6i06IF6K1Qm+rYxn4XPdsl2wdfEklLJ2N2WRRGCNaaFYF+K/+
5uLooJ0av7NrYlz9+otHmP4TCFRto28d+UhF77YCWcs9K7OjLlnBY7aPBO9Q
dm5uu8vNC2zmLHJSeh+2LXrIPEqgArrZaint/mel0om7xNV+zh8X3BfPRQvs
7P9mQs4lkGWkFxg5+Clt7Rm6vJu1HTxGzsyr/g7cTWu1iW1XT/zbXnYQWYrd
M+gvF80+uwoh3D6fnvlOKoSL2iYEskAfD9e0osvmRsHlY10aVqY+99rdC7Rd
Jmho+fSsKKWL4Emw4symgtotBvOz8l3XwisHWkWIMIfBOIzQX6dcc2krezD4
RM7vLFGDLGLDQj+w0i8q9JKm9NzpfL65VyoLoslKJ/8vuOiWtyhwUMP6j/nl
DdwdFrEM6papInRi2VZXmyYTnhxLnS1GwYFa/E3bu4FEXr8+46tQ3rI//Qwx
dpUD4mIhuxKBSzohGeRJgxwdqk5tfUz2GG3747rhFIu1rmvx4UgStoq34yhz
9ob2zBTg1XpFnY07cKuZhZAOwIv4GOiJpOYYHB4IiKsv3AUscAo7DIl5hn7M
z7kV+Orzco2QW7mMa3Nsf+ilgZqZLusMzVZ5YZc+X4/S6aeEwTHXr9nDx4Qy
iXO5b3XfXAcxMa5MllAhRuUN+IkxV06A7vXC63E8g9JsqSw7x/O4vRVmsica
gxxAujosq/559/IBnf5vJNuFiPxCLcLm7+uSNaKRZBdXtQ3MNjDXqdKhv1rO
K6hFoyxcSIcEipQj/EfbovX3kMmBO83nIjPRMpYVJBMtYqRXOoRy9jiQuOIs
qzUgASj7qY53ad0vA29AnlKFeaGP6m9ULe1tkfoqgw3nfsDpEHwP10XGS1lX
65J6Ljn2Khx/L8HDBkrFhM7S8PI1ULCTlBsKNKKMX46uIVxkgKXBmIHnsFsz
EyKwiEjAP7J+IKdD+b+kxpVhOODxxIUEKvL9Lmjgftm/iLFuRxw0Q8NKesJS
Q68F6d3xrlrXoIjEZYitvJrUXQICl4fmh0de6AEr6D4Mqg7CCIJ25LoCIKk1
lU6u2QWXrWTSut6+xNrqy15nPm+gX4g2bdobYtBjoJYCZu1rhGWeAv2YrVYJ
ChomXD6UBZhEHq4FQY2E0zkYJ3WbfCxc3WUGgvk6AtiFcSPvl3gEnMPUqPza
EoOdTPuG8WI0yY1V3D4bGGYVdb6a2Jz1S2uCyAx9hky0jPP7gLDzXgDkULKS
fOUlap4gDEUdJRpo66UudFR0rrnXCywWewZ4kXc5wyqqTfXM9HLaZuFpJCXt
wUAyq3UrHw2vOl3/o9geCXzaIl7M66XRNAlMlhPdrhT3u9Z7C/h/uAYH5d8h
xe/pqxv1tSn1m+5RXu3VpL+HKujkn4N45gjic4HT47dcsNrYeqaTsi04qXJy
WkoeIj7Zq7kO0GsCNqfsC53m+o3+xcnyadOxk8UEjIo+m6oLgcDHRb+c1Ew2
J482Xn4hiLiycoTtY6jF07KhwiC0KFzFARyti/UncD6QxyhfewXaVVwEL2cz
QjU7ADxzOZoIKuAf59baGBc3P1EJaJRV4NtZ3bqzLekiMeecIPDH01MQRNhy
y+qDT0YR3BWYldv5S4KiUME9PzMIHzTPCuxb3+qmBms4WEl1AMvmoHpsPfzn
HOTPzbdDNdwSNem6VHcSUDd22W290NOkpZfR7+h4Et1g9zm8Ekima9Q17Mt6
amTN4Aoii7nuTHC2AMJXcU40CBBa/6T5yxtZ0yWx2aBrkanIoouI7saNLf79
sxD8wtAeeSw+O2SvtPfawPTEiNOrFFwtii+4h04OSKhQU9dISIPOx+LixpSf
pGNU6/Bs9j2DfzDm/1J+SJ10XsZXzqnkSCrBiwX7+YIPJy13cLGIJDjBXdtK
1EfPvxpPjM6s/a1TA0lOMRWltDZWVAerSgrR1XkqGeqpvP0bWbnArkPx8iLS
ly3N0vhqWHQ3xDHOZ72e2lV0+mUuq2Vldlmfu6LLSukXFvXyY3b9a/ufQLK1
RdEMCGtKJJjmeRTQrdAKtzWPo7MPHPoDqz38Ahm8b9Yic1BWFCWDflw2Upnh
kfs8FIkWv1vDeWoWeYNjyJ+8vV4yEHrq2w8zR2YbfdYvu3TMqyxNC+oz1Kuo
4aRskq8yPzyheNZ43NySXKrAukzobR9wj8bDPnO1bXOVlRCdR4yLXiphvBDI
qY0nZixVESsn0gNY+dqVTW6idfKD83fyyLuK/qrpqzBuiN6u80RukfCBfOY5
hvfKl0HhrSBYxKrcGlqXwXTOQ9RDk1kTQRVuY+U6pSlUagz5YLFSpCEErrBb
iom9vSmfUqKuZFmLcwukJ5jO74HwUo2Ymg74lSDXuu2AKXL2HJJrdLx0yhUz
TvVqk9fYUdCAaAXN8ZPf+X3L53A/uMFYHh3zc9+VALSPnpPb7N+Q4m3sWb0X
9mu0wYE4O79Tbpe8gY7tGtwyWCF/DWEe+bp7YaRrXVLT8GBOzYY3gRcw2bOh
Wq3H6usa0FPBsGQaOpWNL1fTqufTMj6xhnsJu4X7yJC65d4Dy40dpiiojrLF
fTyArt5DHFSjb742MjQC6plYrJtIbBwIMT3zugW9Iusv5RoqB6JCwbFFM4YI
if4SvS1Mw82tN75NMjT6aOJKVygkeFMi4EUfEKVJXNflJrlH7yQFWRo7ZoB2
sqpTrdelOB4xFUoicPh5l9L5uA3N4clAFqJZlpQIJYbBHpom3NVdJcaXX5iI
T33jfLBAprH5EumDbuzVAK5SUBZv3dvXHhBjliDPanNxoMtXMCnCjrpECAl6
DuYlx4yj3Bpyy679wZDs0me803FF+WOaw84I5ced95IrdGleefJhBnwbuBAd
YJMpspN1kyxlANiVehHm6T7DJP0JGcJgrd8Q7O47Isaa6eQbtW/MW/IzlEfL
bLgrK3P0MJap6yMsOYcQZeY6PsAVK6qaIUuXLqQ6CFMENYwkNhpFbkgr2x7z
O1S/iLnNlawqBb4UtYdNEoCzcBGcU+HIl/8E7/uhW/53dqlOgwEIVfF9Ka1L
uU2CZDu0sg54dCBePhEIDlWuQBCgI2U2zsK75J9N6ge1i8p0bRulXL+p/eWI
fjqpVb0xcHZqKobfCfrGrwV8JkQQeE8zT4A4xQ98jRhkoyMHu+5HtoRj3ip+
/Gh0/hw1sikT9VTF96m651lHEzcZ5eJJZxlQK2AEp26+Yxk8xmkjmHDvndWR
nXxy+iJzowf6weP1CaK56pyMAIF88W8aHfCrNfERolYEhzmO3FdqrRSg/Bej
HUnWUO1cW6GTnwAnvLBsaF+bYqlQEgad+0ZYLUHG1RTQcnuMXzQ5m1Wz4ToG
I39/tUAdgw1JsMyH6cRzgGXkOZNgegPsa0UWd5XPdNIdOeJad4AGVXGYBwgE
kcUWBMn71wQdwlS+q8MXjwudgvZxrOXkdDsv6BFpeeqHhSDwAI2uFtMfxq0x
K4yg64xQ4ns5VOjxqsA+BF1IKM+cLFfE7yI0KnkBFlnbp9bDHUc8RRFf92XE
a3IZj/aFVzZLDvul3drO8Csw0CaLtlHOBfVbry135zVwNZMSbWFSph/PMBaa
4d9zzjR1y4th3BhHogIi12v7LnKpq16DTHBJeQ2A/aOo2uzEdAF7rHDq+m6Q
s1IbJrRn/ctElHj2dX3wX2xj4S44qUlQTuSLKPP/SxH1ZwtxrnokNS8WworW
a6rYiYFW1DnzVhdqwrkig5qn4EAJWeipN8t4CoVbrhoClZgm2hY1F9J1z9AV
w+U2S3iOLhNeD8NNjXk0itO3r5yPeyyyMxUDDsQZuRqpbYxKUYHvtTBn8M9Y
cK0XgAYlF1IoQ5LBCloMn9cH8gT8gCR8tsHbFcMkYzR17Dqr6jhfOuQ4P8b+
Ix055gHVth/ntUJ6o9pjuIqctUvTkVfFyPa5RXEepVWzKI1zue2uH/wqJxS3
RFO2rVCdt5C+xv9qtCH3KbQD46K4uZn2gQLLlDM6IVxkUckLqAECKlpCrb0H
c2XdJn6B/ORwSRuWhIL9v4v0N+L1SoCbQMqCt5EsyEQ3uHyRn6EV3z3NxX6A
9w4x4jJ2RrNoZBT8jopZOoaPCdt5I8pOZxjkffQYbdHGMKBDLyhg9K2bkBv7
cEQuvCrV0wqNOoby+RE2cpoLpt2JgQxxbMNsZASuYo1BLcicT1tgKsTFeDoa
F0Wnj5PesPXYPQZWwTWGOqi7QegEs6Gn1b947hEUE74kbUGdbEUhAYdseEnB
GyW9UHpv+EuWOD7gJiRv7R8H1x4upIGNiUdz+tbMjes5jm7wmJ6gIHLXHE2/
/QejegZ3fXyX1roRXLwqataL7hx6dFhjONBKvpt2mCgEMj7GSy5xG3x/3KhV
mrhHNiqqTQuNRNqSA2VORkuMOgsgkgA5AEEK84YoWVxHta8GfWc90hdCu8bb
+W5lnuQ0QhbCWCZwJ/mZHBEUIIgaGklM0OspztkMw9v7czTgNBjLyUWpJMmD
eO7TMIakeVhO6vSCHIX7EA68jOjmWmLmZgZ05aISNsTyjUwoW1lUgze4mmPt
tNcsaS/iBpgAQtsI2i9PHQl8aCeWEgquMa0DitP9D87Y7GoS2grZvIeI9WUk
TJiMuiODw0yQN7mz2EEIzNVDMplBt8FIf+NlSOaQvOfflXAvTIXV1ZjEULPG
47zqwA2LEI6iQXbeH9HxKGkVqN+MgIkPY/TvAFw2Rue3P1VKuIb3tbgaLTGJ
P0fx8rv67F6cQE1OhvaRb7dUTNcCCgM6H/X1wALZ+lOGk/Vf+9GbmkYKvgWF
b176IpMOk0F2Xy4bVtn582wxmw8b5yYENzVZsFmgt8I/C4w/Iha1O80Bn0Ic
H14IvlQz+zJBcIZMHsmOzqhMu0dYizoU68snSjMiHxkEgw9AgSQs47rUGkpY
Qkbdpe/iqRl42ITddz7YVc7tL03ry3U68kUqJAtvY0LNmiBUoKfZgXBoxPRD
UfHtITfsPZh71vDK/kuDmdRVopCrzleJU8V/PD6+OEofcXg+24xgndn2R0HX
AIomLb6YmQPMEBHCdybCLHgVXP2YibsnODQijfLgFiID3LTux23WGGA5s3Ye
aGic8UA9eT+EUemmuFSyT2ieqoZfo5FhKJ6JwZ5sTSYPHDGaVNtdS6eizSd8
Fioiazz6vaeVn7k66GfzR1wQJsA+lhl6TdBPvz3Bj2y9POGaRmoAZ/BUAWAb
+FA6Pwp1jrZvjyWuDFfSCT0SIGW95nBASHj9QX7ci1jMuG2O0KWFdDHzZ5oy
0C2dRGcsInMkNJnySu0EJKN1oGGrrobiXbrWYOJ7OL7bIChP1Bbn4i8k416U
RR7alji+MfHx0fdj92xvyvbAXeNIOxPHVTk/WEe9npn0UfklbwBjeaT5d+pA
UnsCkMZG8Tc6efPURvI0TDKOnSCHvyKJvDc6QPG1JfJ91W7ET0WbXeFsgiq+
QEiSxiQKpGGZutM128JJgJ0zM5q7k0k4h2kg/QoHe4/0HYTUe2tviRCGxhff
Kb/4Kur+YNnrcRwIXJotfb05Igx3gBJeRfy4MiN3G6Hec2KcdKpKa5WHMRZJ
JJaHMlgt72/Ls28us721pora3sBr94TQ/9FmZHTbCrwO2skRqeJaaQ+Frs/7
qDbStUkYLqHRAhvgWGa1aHdxVT26YCW/ckWWK1+BCkfdp/L5GnPHxwGBbgv0
bnLcqlkyVMSZjQL03Bj18937MEV6bTN7TWIc4nqQ8MldB287GsUbhhHGHaqB
OfQcyASElrW3kf2yoqEtAddMpBD1zQ6sIYWMl8ajDZcCZU01+meZR1ZO8IcY
CvjaWjiEZeYs4PmAp4nBa3DReZlI1bq3f/UIW44k43Wml6fVS6FEN7m9Fmaa
6WouxKZPGAmNHK25s1E6ZW2HlLNlCOlUTaqc3NEvmSA9hDFzgeqPmLhjmuTZ
0XgKS1uQTwNwdYVy5oe1iTyW5+4d9FdSwDBUih2hVMQRl/Hvpk0r+tAaMdSs
lC4e3jjMKFvYxCGd4FlksON8N6shCdP9vawBO5HiAkBd9jcY677FrM9TQf0Q
cf6hxZKmhzeQzEHeUoS3bu8FDomboW83KAB90HkXSRUsr2ImmDSkxQi53Aqg
vOP56xGbjcq/u1busccyrmI7rXKUt5Nw//F8O51ijvLZJCiQyXLyJwiVhqYd
j1XUQ3qrY1+eK43VH6IEDL3SBkiBvsCefianKQSDhc+ThX1Dr1VJNSQjxQJt
n+amE9ryjjRYKOeuh+myowMJplce5Ju++lZvVv8xC2a2xE8K1RvasTiL3HSv
K7ctsXlG4VbQuv0p/KBolzZU/flg93x1uN1N33xIcWTBeymWwUCkpmUuhrbS
Yos7gnt4saDrwQrTNKcCSUSkfdG14ZzmvvWhufz2kRA1l8M/clvXWZZerhUv
EsWjOASWETYasFTc7jdS9c56Pff70021z87qyY41Cg/28lKny45ntmkGfNX/
eMB+uyX5A64o2epFKNIZCp07lWKL46OEIdvPTNTYXcouSuOWfk0yz4OcWfgz
N3fs21MUqpbhv7RiblwLikIGdRRkJt9ORpG9UDaAjSwz8B8AVFJ5/o6DL/cA
84U27MFvmgOpMR0XU/Gqoj665xmqhyU3WSQnD5AWYV1iCrXA37S499rigASe
KzolkyhGSoW7mNS78eoflYzU81MJS6zdr6AOFdpBYS8mPILeZncDURrlzVYF
wauiwtZQz2N3iDsN5Jm3Rjkym88bZce2qd3dBZbYIJ0w8DqqRYW1XWUZVA8z
9e0bxV/i2rd3l2c+Bmej1cXspjVil5BdbgN2i50DYFgiVLNX/0FEE/BBR6ed
iB/J2ZUyWkuJbALJheRdN2TgXYuOy+oGPxTZaUoJXbiOrK5i2W8PDD/jITL+
4xYQNkupRngmVfudyCU7fTXGTWbSJHhbPa2kMQM9wyFjR/hTEv3dbQ1m5kvh
xY3vJ+4iL4lNX+ZA/fPA2zah6Cct6Guw2U/WDfTcaVSwMq2KNLUbrD6BfvED
ZOQ0cesnSF6+Obn+8oXBDs1T65QMJrCqvoqF1SpEp9vbcczhrSPex+C0sMG8
uxhz0P5CV19C3gjmcmYIuaEV+hOr1nPNy+4mb2xt0/3LXPeIwhr5JePjJw3L
gx11qKA2XrseOsaIq0F9tuAf53mfT6t5XrcjzRK81N/tni91AEbmh7kGXJk7
XaFpdCW4ll2nOH79E7CpFkhbcInkZV12u9rJR/uPYT3viS2YtcL5twCLsRUh
pCGRbzk16JXtKl1j4L+1+mmWMT3sI75yf3YGy5sUKogs49ay8E2bxwjk9MVp
6b9Z6VSg0twlKE2DACsPPHZBJlI8MOTIPbRVcU1cGcMScsHcaNov8XDEj76w
XD2qHy8S0bAmIqL6a2fXlcXOQ2EqBL4dKfj+rQ3rdqmusCZ30UnKUmtNREoH
BNQYmMEsH6AmuR1oXIF3fyyZHGkjcm6NHaPo3+KyUrM+gUbTK50fWkBIV321
vxHZoV9TT1fMFDAV0v2mwYZzHVsTIlLL0nYSJyYjqd3+kIV4Cmt2cgvBHaGn
E4fowi/U3dY318W9n3mlUIY4EOkzwLCuuPAgQ/geo9Srwa18n/Tz2LNdeOQ8
jSZvHPiESOZL6md0Hzg5kO68XIxl1ZN574t6kcEaxfcPqi6kwhb/EHSV2xmy
fWvpnWjNC1Xb8lKqCZ3leg1QOe9MMhdtiBs82TUmWbWNAIbxdC2TWlCCsK3U
/42vKf26T8wb0Q57BcPpB+j7w/T9GHxel2Q2LqUjMnBNhZsm5kr9JW8c7I61
vY9GJT+1ZEOpu08+kHsiBrrMzcTy7Ou8bwObgNgA9m4PG4NIhaUlYxrMX+Ri
9c5KP/s0J15nkVRzGlLTas9/qOzS3/ZDYy/wmdNZPK46DVBHi7uBNgnuLGfT
/uNvM87/gVCEWhJp6wxE2dt944NlrrMefQ6YZDfVuQp77W1DZXsMX9deHYTr
NYnpzVC3/EYeD1hofQGrvt9bNOfD4vqBAOGipwnFE4XIS51grg8rzp+HZu1U
2aU0DKsu/MaOr1/O0Z+NZrseDAzCxu3jiLPnnx7IKFobYzqFrTXOriNJgKNA
jqt70uBrhWUAAA9eUb9TDbT9oDX89WoB9+2k8b18xSkU8RCO3WywxDXqh9hr
141BDDVf2DKNqp89UTagbyMPcTcAI/PLsGxvHRpG6YlzIKMcp8OiBa3sK8hc
gBeFhRuHKIXV3aB4unp3sJ7qhKi2lMgOoS8ZoW5YGwm7w+ESjaQHNQJdQGXF
4W8rJzKGhQcrra1GHmbx80qEI5bPLv5Tq/+ImIFE8yLae+ZTbTHXV1wI87bl
Ss3U253LPyeQOocLErtboSO0X69bzQeGNOTA6Uoa0v0/s05tsDJ0gok+l9E0
PXyYhESXawNSo6UxqRV3D86BclRs+GirMWIIG2NssBmxVfBj1MNizftSM/7H
QXvzbd7l/hhKx4aRAC/O3z9mNHBbJkV9+c2PRuRknTa2FY/e7zTZncP/C+ua
LiRVGmOlSOT4cheQAm34XB7rn3i72OG1KOF+S3l6+gjCR6g6zB6Nwpmn40Hc
0cBhZ8ic8YChrhiNPsUypsd8ESBYtvRRN5m8guj0XBTdnALme7nlpRScJFl9
1q4pvvkGx4AX5Dy2Vh5GSj4a6MME6jjmfm00iWf/bZDcbppUffjO9eiRzQBa
ZZbUfCCMIdFxqOiZdi8RlppMTFltjvh6XCzn4weg7L8aE6c3wDytYcPcE/4s
pSLaH3oK3OdkXZIFuAMn0EGprRClTygO6SC1p3y8c5xT3ycjTW0MMpN41jHR
fnJDzbIovo9x+bqpni8b/Y1cpiJmpHUc3eDUWIBva0m1vhVoYSpmh+/tsL/H
OIG7Kad1e8qgTVJ1xiiw/V/hG7VEY3qZ9qg74HgPRyPE/mkF6+fAvt3my8By
v6Mj2wmkHzI1b1aD76xAWDWg5mBZTbqshTa2jVciWeg+FKUwOUn8Xw3bo2cQ
+wvxMmpFFJes+kFkB5woV2a1nod3I8/7aePXuMCNdLVS6KqeuS1NwqwlxQra
WtMweJJd9mTtPsW+cafWrlKfGRl8/v6Goe4zqnUbwmMpX4988rMNFEx8inzT
1BG3z2MUhTjPDrBv7Z7wiHBzg9PY+avUP5vkqrA11EHqkafMy6lsk/Zr7woe
K9QQWEiTnVaXlQmFJl6gbLZXZbTd5mmudxraxihjA616P/WUn921QJd0f8K2
tC5na9FhHuz7unEeSAcIVZDT8DXi8njuP1LMXNtpP/lrfNPMs6/axk7k2H/d
XhNlu5L4vxg3a1Zg+GeqvuGHmmZeJ8Ah5oHQ4HB0U9i+oywhnOehiqQ8e/gK
qkUnIMuEy66pUreCYAQQSnVc9lvhrjiQT8E16MjUl+i/OzoUPmztgewdagxb
hwT8pPw9B2XFMy9hQFojyOcgOa0WroswsRkW3lLgGfvTkVgYl+FQP0Hrv4xK
hAu9FVQUnHSqtZuPCLIvtZ6uvB/RmyXe3CqS8I5aCPoFMgzvMxnnUe8VTvBs
6gqCgHJwLS9LDlFwlrc0fImQkcYBxh7a6r9PrCOyogIYSU4+4zS24iqXkpac
p28V9RY3cMtC9sixPX3IbsKTeWbNyDJ4wXijZJwarhCidluYZaCV9icv7bCT
xZ8/JbOY0CnrAX/O27hhrmQYCYP3HlzDTcGE+S5Upbc4g+PGHK/nDCjzeWSg
Y8KB4/4skRWO7YNucD7RgQjkVwI4L9f+eff06jj98wm1laSiyUi2pF3QIyu8
WBUtjGAvcb8OTj9aqwQuiod2NswOHWLa7V/zYaIOAOgt4YREmcmdvY3Ipbow
1lsFP2cbj5Q6POL48wALjLGh/LKWsCW6pISZBMZggkCg5dAoN+kWWiNcihTD
XtkkMrlA9fv+ZuY1egw/0Xh1gpCKCCBKVmiPxvwSyAxBh0vC+aWoZW1wEjl+
rIqrb1BpHsKjs8ay1zYnmTr5whzyn2csJs9LKpFAgpnco7JoQjaMYxV7JLB4
cJiI1n6+0hdNt7mm5gKpTgyrGCc+z6GY8VpaufiAxNi2iGoo8FbemmDkWQOj
hTT6HOr7e2w7+Mrqrogv6av8kYGC1dfJ1el7lxCvdvzfdakCynjiwG7qII/U
kgwqkINpAnng3DNnvxCUKNV5XJuGF4haWFCCGz6i01GQgSq++OV6P/N87YOz
hXiivzWNtySd/FoHHWVhdhjww8AfHsJhuM0/K4VSSrItXm5nsNLm1fn1U5F3
widhF1w4GRVrpfxUu16R4NkoYOKEgYr/i86v36qug1uey/wcIwHUVaSjnroh
SdGC5r1A+fDyHXaXPbbwO6j08uMl9nxU04p80gBJevH38aJOysda5Mi87gM9
9mmiDrv9GKkQuEWJSYY/lqmOcrAqiacOHPtuMkWMbXVA3U9M7lixRd/nd8AK
tk2YVLjIUo144C38yxDkJpvA7H6CkkZAioVBWWYcyGVxRgk9sXfJOLgJhwjH
LaZbMzuLGWhajD1InfH6PwgWx10ZufSwtEI3HQ5ljAkM2HelQGIguvduBX4j
j8E2Q3NlHOfnsYq5K9si3XPPQoB66/fTHJHmZOjiXNfimsFK8nrRQRdx26d1
HMaQQUh1upOlY9iDyeehS6kUjcD+310rL0H5CRMcns/7zEuwgrKpMdm6Zvqc
eeAn6yYxgYgvx/SQvMYvVnx3BqcEi0jCPUOrobYdZaWkHFFRmm2U/ixKYisW
VPKFL7Bm6GKLFhfeB40hWVuBpkwvNo1yX1oOQ8znfGDKd4H4onRENO3fJ3V3
j8BfaPZqK2fv4Zm2OnoSrGUlQgLo4Ldf8B+ARf0w08aSVcV7g7IjeJqQjM5d
FqBMyVZDN8q7Cyp8IdnhgdznX/8OX4wzLACPSxv7vZzMJEEd1to5l7pD0Pim
wfjtKOqlr/i5UJiXf16UR6aVhgl37NAEfnGsKE6IA43QQ3svXBqe4AbiBSFX
T09YVOcKYrqAAI1zQ8lvybN7IOIVhyjd08syr/13oYv7X2+u4M7lvHrnR4NC
CiL954PZL/v/nKocwVPSRO9sFhW/sYEY8u6J9ajH40EOsVwJ/S2+p7pstKzB
Tta+uaAs+zTUTLd5w68VuRLC6oP3dL3sJ4zljEjsY7UBprlhKYyPF7B6LwMJ
Tn9c3Z4K8K3xbQPDUddJwziPzN3EgRNBdCJZH77ZaztpHP4b3JM48HxbHlgT
C3z5IFGiokpNSETktOIbwk6ozR1LioZOWKfQm5skt/SzXWQ27Ey+FuO7taLj
zErLrgMyAyZ0lsmMQVHew9VjEuw9ERRflnTkkrrFd1gJjSvjbe320WuuBMBa
GaTHQyt23sV0M/hf6GJsRwjLOR2G/U6zzJRLMgwWGyH54fh7Hg03dvkdOi/L
IfPMpqasjoY7j/0G6MO0+NfOeGpcLgEEW/k3zBN6IPakGMZ66M9sbes/0n9D
PwlsEvdQxZD2JQcDPQdxz/EjCCOTPgHa+ag71AsU110i+kbwazhvKByUgDg0
pMoZ4livEZjMrZS/RZ5e3fGkREmuhG5fm/V0ZSVZUfDFY+4UZQrhQX4wh+0u
NsxsKykznq2ujTY/TFAoQglibiLobndxVSLYxzl7IEUZnzGaYSEVFwmUNQp3
mrGYYIUUqk6p9AhWoXbn9sT/XXTxvzXpIH9R0fpXL+O+0YFE01gxJFAullat
oVtPn0wSTWKOvnsI2pDFohVlfWcSMcnglscS5Cv9Us36L/+oJQazJV72nNje
pTf3OuML498zH+DChBQPVTVIpPqqZBrbJGDAgXCatj2FZ77T6jmf1UmIVydb
jEW/i3iDP403a0q+LsuwWIlG9pfVu/kZAmDOP8XKi+BxC2e8NV7ffDm4yiYD
Ow9KHwgOUyBVuZ64DJXTDs5cGrrxZa1oZ+nBbVA0WKNodWAdpIy53PnQCrZf
ZqTwEq2EZUo222El9gKRyX/F8yfhPj4vzta5+QshhcmWiYJ633CDR+9ZuPWv
4odd7WO16yJjhltagmimwua+EU/Nc87paoHFuRAIUmSJZyiehmOOxkwai+No
Q6izVcaS0plJlppCXiy3rY9olWB5ea0w3jRl062+195JbmLh2D1oxMy4BxgZ
bDDgPFcq00t704dhSKo/HSq3lbz4B5fBwsgsie2/6XjMiuoAM3HJfCvn3pP5
LmJIpgJbFd/e1NuAH25fnndWD13LmrK75qk26VjkTaK1VipqTVV89i8mHknv
sigOPrclPj0ZmgwykPDgrJ24mJMtwEyuOrKPpqp0v62eJnNO/zcmu/HTWvc4
cmWcWVuXjxExVwFzvq2X4qLK/AZX0DktdF9ZvkkG8oI/84rtOVgMMtdnaysH
TUTnnlIBCTfpP4YSqc9XTyb5efiquNaogU9p1VgRDVRkZgUgI7OpSdZL90Cq
XimVlywxyE9mnL3iruHlgD8kKNvtyMXmG0L28K00Y4e61PXfNEJNbaGqimbs
AOHXLyxNOpJfEiS2TEkH1scwQLm3/J0bfqZ134o0TExg05UJTmQjiCGxCUBW
dtyj2rFqYGZFcuVrlxeePM2Ku2G9JOkOCRgoXjJr3oNANeUXdTAl9qqNofbW
kZPvgOzDPhdxUXa1b7bO2JvbPP/xZQnEohCov7qjAYplX2n+zQJoUu01xPPf
ivAYFiHScQ8OulbnwLxroZRM70Bzd5wVNso8LVOCAYaCqefUUeEnxTJCgWw2
4l2q3X0RsbaMMx/tX2ZjN1tZLkfNeIaaqvwDpm8p7fq0BX86+gNuT8SAwpIV
XdQnOq0Msp3EXUJMPlOpRyST/weN/+/5m+qcka2hUSP8pCh2xJbZr4DnASaG
8BDk8df0T/dW85zU+VZNiSL6qAVwqj8k9UZk7MAm95IyHXZLZ9NbSDkx2XOl
UtHAFDMj6k7fn8Fs+rYbe/yyfVc+yX9oqIUoALcPrEmx0mAV5eHudJPEyXBT
s6rsxtGB2R6GB06ar1ix/MSn5JKu3EpWME58ysQYBmUq80crSPF0TVfD/QxW
F8j6mM6miM/gyDqXX1lqqj3UrlR7tldlHprNDQmSCZkE5P102ZHT/FCQ/nBK
DLifnT6LZC196wRztbaOmW6BihicwZvftyEnkSm8KDCKN4stqaRv98SvdgyF
IhCbY5N6Q06iR3HJFvEwk0ZjYp5SM/c8qCr3IDDcXOLcjE+ckSvI49OHp6sO
3XzZ4qGtnjaCSzd2/o82NvtZtzLOylIm34+MT6liri0FmLRRCsa84XmAYaRa
/AKdVhKr99gZp3ur0yOnug0ovuEsiwALf6eB95yfBug/ibSrjY5j63D+LaXm
UR7vRyj3E3j6zAqJ8+aUD5JFhPDXjQPxLDj1kkKe7xqYZIQZQ8wqspdHC4BV
QccMb1hr76g3/ZAyBnQNghiGRQHsV/LhKjyRSfFhvXHFCZNDfT2hxww2J1cb
Od1pGwR1nDp+dpklomvqb1UPjQzA4mNR3CvXcprOP7eZ+ZZia9P3QaEi6yDZ
CRaMS2Mt6LUkLuvjMrnxhBOSp3mgrsddBODvaM/NGdhUeZIeErox5Y0I7HaI
Pofvt+FQ4wf/oNpV4p0g13oEibATKJtSFlsIzhn7ZsLYU1hH64K1uBXDmc77
/VHjrT4jRxtUCK6jE8TXEfKQBXJNeJGrsQ8y5tPuUefAR7xb8ynKYmQ87gfJ
r2avSM6FoXdp2WwCeqt+vwp0tZMHrMj2xOjyI7yZJ4bXOl/UsosRxQ4LbD0g
XDv+q0co46CeG0/0a8U//fA/Ep+DYvN2RQHN13lRepXOcf9jqamj02ggC9qJ
FVWeai97Vk7vKj+5emiflrUh8zzTeFySD5/7+I/9nKRFkZgOMe3I9FCk6hU0
DupJbU5QCP+8MF1t5YYvGkbvimOh3PX3GJjCx6N2r8uefYwvWfG54Vhjadhy
X7I4CmiFipI+WTgSnZyAfm2rtq31IH80NAoyE/BpLOtXApGDdHhBpojpwhPn
LWQi5CvvJaLFUgI65MKqWAh4KNQKIRM2BRu3guS2IjogSc4FwgyqlgAz4qyy
mbC2ANSszR9B13qIJIAUGD/Uhc8qYgrR5tTvz9S7wqll+MOpZFwvBxKn0lg0
4H+5Qp50PDiAg3u9qw9LPiuavkVJIU5clWBWVmVqU4zh/SgngPn8jWEM9Lq/
z0XjaD6npJ8K97FaSIMRxA5D2rQnki7+b4NRLyPpIf2oM89V/cGicXCjao1W
Ff2GGBtSjRAOoyJJCtld9TLfcy+p1jq2pzJr1ppmyPOMBTU7xBNJ7+dhlB29
Py0fcu0CdwqMo7pjUS5EL1zztfK0zdqMwy2k/+GLJ2jUoJr42S+nXlLCIlGU
1hMehDNa9TiIDlXpuAax70fpc0uex7KrYFUd35FfPLTNHwJSIBLFKedRDKtq
repblXUidIloIW+qMh7deqN2ea+lpyKCRY2WPY3RWs+HhSu7b3iVsckQGxgE
ZpKbIFj5NBCrD5y8kLlsIpN+OJLYQT/vRTQUQlY1wFJgDSJjOfcfmfG7q18G
mRpC+g2uJoTJnp+fRkm8LQDNZ5zxbUm4DgswPjWRTm+n9X+rwyYKmz6TCTt0
/S2KWwhbl4yUlNABJLQfe9KBv95oloHaOu7GWZAGJMHfQQU88Axc81LCOxju
P43DTqZ02EcfQI1ii84WKfNjKwkxkz6LCEXZ8CLak8F1SXX14UKdLXn/Chx3
dMTJKFvtwH8QhXoicy7zyFLZ0vdzvr1hGLoFMIIyQkje0YsbRhqXljf0jSFY
9X4VlAcmu7lCpEPZ82/y58gPQZX/0SjY/IyKR9Mq+sZvq0Cy9deQWwqMFJzZ
S+bmKy0RdcC3vgWIOMd/pw1ydhcx/AV+LPgQ16rrM1R8XdwtENDNVB1Zf3W6
8bLY9cK8lZvkGGzdJ9C8xDf0TkM7KKdyVzATsv33lAJaa7K1J6UwuKkcNjHD
CyMqNchs7J3cR0ygJu7eiOjlM+reT43Fgkp7WH1WqwxlEfEgt3bKB+4QgtcF
qmSbmvTExxHHSLCsCLOmXsh+nDGNL7ul1yhIh193usaoJ+IKGn2RL9o77hjd
pSXuv/1OJhqgVirkQeF6l8Bt1QspQb7ZNhEkH7m/67lw1lxtUSZj+Rty+Ezd
2W33awIYEHbMKa6XK0C03oBbjaHchmJWMuhxXjM81Qe4Cq9ju18idKLH/xQY
uTbuyoB/rfY8x1RkXoIauGny2UtpoHyiPS2PPUAQw3lfadhGRxMpOifbfa1s
52VZYfKvqbhkWOYU3JVW10NNwKFc25SKxGEhboCYPJHJHYvOQjbgq5ohndm/
UuI/jCgzkYGCMuFGNanlng62gbygTaqKmy4nJjFnnzWjVKP/VHvYTLetu17C
1xipi3smgpcrLSb6yvux+LdmtMDioBxebZgOrLi0tr52mgrkyj1+yENE7Yo2
d/Y8ebb6DkByHPW3sdyRt70JrP2oS4QsKgQ1Hiz9s8YYvJxBhomqKOnBJ/D0
B9XmPQaDVWJjJzruDdHm+6QxooIFkAb1JT3AFpa/Ry2MaCk3k7osxnPoWm7C
axDJe0pN0aJ84I16mQ+XPn+3C5THZGAS4+fa2hJocEJiqQwnnnJUw4Fo0WLO
xDpH8xlKpwXHE0/Nk58KMC8JE57ZXtG3vVV5I5qUGIGtHd6vDLiYFLmYPYqO
/VRrUg4PHrDC9tsgiIGB3USUDumSj1r076V3JPECzlOh3iPc4YXqKSysAi8b
2zUY6eDBPLnQDKVEjcKbMwuu6qy50/EwuWyaod8jUljTHEu6XYnf4gySuao+
OO2jz01Y1e/E6ilVIlElMgWWi7ZTzsonDadMVIZ1Kfr8Rx7VU0Xc/cont2dP
JF61pXMCMF3YVXqndQpwgQbPyA7nZhO1QhAVQ2npiQ4twID4l86lYpKdOtcj
i6BX2R85md+y9YPw79d0rB2BPSeNcA/RK7CZY+/ZOj8N7OKauKaL2l2kSfy1
GmeXeP3q4/wDC52aLnbAMbmITCiDjTfBL8XEnJhRBY+TrSHWkM9O/FbTAyWC
yMS/ZitV19EQUDUWp0y3hjcNIYJQmIerbfoSOen5OrOh80OrinC6jY864LtV
qWweDummA1xtLxDaJj1OJEbyiOg/bopN4PSb1oKZP1d2gMhfnZiTJkULNqqZ
xAq4m1quNqQKKcvN8k21v74/ZyvfuBBhTNX8u+Sntm/5D8ciRFeVTnHv/0sI
5S0BPfLxTo4xNGJ+0n0Pfgz1/WAblFuHJk+CqiBZ0BVdj+CRfKYQ9Xlvw4yS
m0Uujll7WXQCttPk9bNUCfDxLF/FdklEdmmT6Gi0VNWCfb0o1DHEBOdgyeKr
LOgacZz0TlBTgkQ+kqWHu7UL/XND9jlX7swy+dXkSs2VH7wMzVevJIfuSHyL
BN/+SsjfHb895eSn6QHJ3LMmde+cY0xvIrAO415MpSuHQWOElqpCBh76l7d4
aHVK3HVQ/W5nFw2itFUFihMEf006NIgwaChRjBVZUnCIZUZYTFOKnjA/OT/M
j6lnMfDrWkMkHgRe5NHv7G06cAE3YBijhqX6wxA69wS/Yo8N2SHL6BuB4Adv
xONX6LVT9MeKnZFcWhPpE62Aq+yQ/FrF4Og1eRB/RcMCtNzuaTd0dzRpx6th
+u0ibaBV/Ll7/Uinc8jxRCW/FYYbp63bUJZ0EfzdS7iDyI8P3WJ0k5OpI5fp
tnIh3+ImSIbj+zHTiKZcbLlGbAruSZEIQrr9gUvGwYn3YASYiITVytMF0eJn
G5PGBmyE+1wEcX8ujLnoJJOZlawQPwh7GlkbG/XSbBglDgQf/EGfVg+MwLta
KY+s3s1Z3QgjtKXtfdbheGqv+UytPK4XWsV1PTJ/t32YJrn70y31oi3Q3qm0
77mir/b8t2SsfH976PvXgECH9k7hJC6zd4SiR51UVQBLBLzCZatllTySQSkq
u+O24N2OCttiUwMV5MYAo0nj8DX0dUmI7tlwAsesZmFC/gO/B6YF6A5f9qIS
sZ7Ombnh+TvudaTniMvEBPq/G5da7HDJIFJGZspQEOupVltoL7WFXL9sMHf0
QLbWQEwWYUx1dCyzO+GRy9jVTvC2wtI++g5IGX7lvCsVwbU1Kkqhd+Mzm4Ew
LfuEfHrGKSv2GjWGuzgKq3uR6O1BfIXw1p5dATkMBok1dMLQSd0JL8Qbj83X
XZt3UAPBU+GTUPHG1CsSDDvgqxDlmFusgjFD9eAaqMMOVOqXzVD1xbcdbyVn
fhsBMtq9dSnD4EjeC7dBQkao2VFrH6/OTqXVyYmVF8B7lW9E+Eo847VabKDh
8BfSWYKDS4d6Rf8rbYQSdNaM+CTi/6mm0yY9C1ixDFS0LDyssePoBDvoUBgo
wGLGxbeyGq1voHQjKwdpscC04HlXpzxILp9o3bG4ODAHTgnefbpy/oQ+ElAB
NaZmzMqOKJwNxMbvgWQmrV/Mm64aYeCLt4lVJZB5L6GcwGrY4c5Vy1M4wVG4
M1Z3XDD9WrBPnlD4gDHyzyMNe9vpqgjENV9nTNaHlE7tTpeh5lxBDckwHSMk
F9dTSzNacq5ILWsgaphFOj6hPQZTnaz932D61StsdomktQcmTOpJQjRM6v1u
PGzgA+IvXJ/dUWze1XqgzIVqKsX7xxGIhz/fRuUrJd/TAWepohJw3Q5qmNRy
GFm6oRHWPYPijUDaL0Wkdu919EDLYxjsZTFaEBXUEeoDEpdJLb+YOLs9+7Nl
bUExn6k+uyXnw63yUb4yn3nDcG51qibASxCamkzln+pSvt/OH67ofkCaucns
GfHIGHfTNinoZjf/ONJXomku1GZdNbtQ1uCbBiXLG7IelXG4qoVqLVB2Kb98
cXjDwDi7VXLiWovv++RRxMZheoT93lmqcH7cPsqyoMxWA/3rwaMXjSJKXgu2
n7/7dFBMPSYwUbNZqs9cFUyNO7d7SPcgZHw3gnKoc3KQKROo5l2EEf4r8m3U
v2Bz+fVlp3hNaV/zXp3smNus3zZJzkrgbsMsT3OTlw58V9Lu9WBiVxSb+fZf
wXf3fT33ineRobNSBkLp1N2LwRAMqfsxpfaBe8vYgpqacMm0p1or5/p4hHZB
2yx8JKzGmyOuQGJx+QVfNgW83xdjLWz+cRoCWMnSl2mMgSoXjCNHDBfQdGIm
4fYqNR/T1SqfxOB1lJ6Yb+JTupnzeVQRWOLWW4AzyqR2X9RnD51jBFR8qx79
qAEXbzXIiA2G+rco0To1UQM8l1Bv4m4Cfd+b19wybmYeANWzFDq9gexs/Te3
PNGWMZfHDDYHk09PLC9MBeYqHKRZDyH88yxnFOEK9bLnivlO2iNXlfHr9N0x
yaNiE+7+sg68ZapXWfB7RBY09S+D2y6gavo+iuJZjAtRpn0yFymYtz/i2jG/
j2AqcAKA0ft3Og/upC6qWCHmPGIwwyr4fS45xgHzqFoPy1KjjU9Xy/E9P5lZ
PGM6TNQkIfcOj34t98VzO0a4e+6z/UF0rmRW3uURZDckfiDoKdwHclaEvb5c
PFKU9AtndbrUYzcG+Z0k2Y44qzwJlmOR14qGFe8RmDY4oTojR2QK7MM5K3Z/
BneQyh85EAQpz+AsvyvtUOQBEXYXaXECid7g+5wDuTuH6YfnxygqKzxE4LZX
1+8eHMP5PbXxUpVBzd8qWVY09PjlU4tMkG3fiD3vnbsLNL7sSxKvK1u/L0P2
Ac8GzE11oeWIdCdxQnCb2AmqlArtxf41MaoRAv7JUAwOEwSEiWgqUi36hJMW
SulHjkB8BPzjalIPXhGT9g5fZIqjsGvi2Z4dz426m8F8i3Ls0JXdSQJz7X22
TsEiK4/3s0sYR2lkjPeu3aj7wGTEImUtIs4IdSlWeMVVSEAl3/Ss1yRTRQT+
bf3FcLcpCgS6kEqnlFUGfTgFDWHOFfz9vJDALzna9Nu+DZ8UQQCu+rlZqECb
eGY/dF3tPjxO2cacee+5yNFek2iepvPAB3vZHdfj84Wv/C6sjves6YypznJZ
+ilYbHyIKaVCec26KmTezqNgdENGn54Ro22gHqYEqVBc7ZHw2IDKcLJIhSV0
kBJde3xa+smkrm+8qfNNrWjgLYp6KtavMlnAAe5VeEIzwwk+hPCV250Vn0WV
E1jDdtd7M+YhVUN4WLQmvYVv9P0jNoBCqt8ysc6d+Lju0iGrRCj4SD0HTkot
5NJW5STCoO8pxCF7RBD9qAK5GRnbyqC1I7HAHyJVCJEk9NSrqTO5hQnTTKkN
Uri2lTHYh+//DpVqrKn4YgLHxMmhxmxCNvyb+9+BZbhgLG8nUBXWpra8//Cz
pkNPh892GDb7Bq2neKTL1iAY4Fd0Xwugk1PW7fw1zBp5n1cAo29je2Dpi0ZN
Lj83ZAD2zKhtVlVVPDkazv2SND9ZxfQVRDz/LuxBasmgeg/SlSsi5QRLVjHc
Z1hgP+Tyw1uijtsd4UPI7vbLFslX0akx3MZ83i53Ryj8ZSQN7wvMAYOE9RPX
tpQqIreHU7CZlFmlvfrXLJ8pYAq2mPTXPFmM6uFJHIFZk3Z6EECl2r5snS86
vilBbKx54+KZTtDv26ueXwsGYQlSgJ9ufxNOyGZPdWkHuIZugT/7nX9qgjlF
ESi2Va7xocuYVOXhpZE6QA4yMLf9zCVVZwD0qlPlPICKr58FqUagpZQ4569u
h8CWyOW7n2xvJ7+RkeFR4HDBZdA2OIIDQoHgjJKR6+7io5QVPo87U83ya7Hl
YFPp303HSWxMnd3o/HnzQizM/JIIAw1VyTi1dnBjNAaywLnMsOjWrKX4qAy0
3yaFk6v7BMhbUvhUEB4tdGus0eXlX32PbtyEPbTiU4zciWP9EL+DfdQA4Knw
244ZrWagp75g8/+H1szOKKNA+LRD1mPGRma+w0IPQdjPBPTsI5ONci7qFBfs
rdZhRhikSTjNpRxhbr5ArTZ9aPgMe9juqbliMssVbDVsbLfvMifTeQm00yh6
/KTsoc3wbUjbmT9jUUx56tvUMh1TyNI79hFvKvusXAu6N5iuulPMbLUgw3/H
EbMfFLN9lWldQLuRWlmCTlyNYku+nE7gutXzxh5DeRedWU/hLX8wWfVgQL0d
m0aNhF6034Ce/BFT33xadGnPg6T7NG0fS47umDMnBYu6MjJmYviRUfa7wyLQ
Ih3oU+SFqmtg47hfCi9dzQ6gWhwbeyYVnvIwgrSTTKfKwRozrMgi0wxekLZz
JJfmxUovPR6YKMu4fa7mOl2wYphmioFtYDQz/b78vExNPHfj6l1mCWxhGMab
6yY2LJ2kkHf7Aq+wDcNpiOaPkHmseM8eTuT0J9NEiMFryoyThhAJ6hDKKZ5M
p4B53R277vKZCj+9GE4mwH8pmzYtkkHqn6T1lHkgRxyFDzmHpCGR4fLtC0qv
7YRjXWOxuRYvwlDWNutucGbjKZiBkfAJK2EZtAk2hr7FdXMdjVfnNF9/LYW3
BfFaiTkSoKE1CfChsXpXD02DKsmQlWSxhJBCJEoO4hJyYkLCKqAsIy1Z9YW0
OS4fTCiHcKy5T2rj2T2eQg453b330j4jakgealoeO2eSp1oilvoPeMIr6DA1
JVmBc3Im6JEWeNaYJ4k3NodLWBJQyxB7FITGDRxWX7npsmMHzcH5jIz6kZwj
lil0LomXOypgjUB896OP6EV2+OJNEzdOG8XjnU41AO1qnqpvzHOdwx8OhAxE
KEB7T8ZG/CFN8KEBe16w7WMwlWOuGbdhoSHs0GEkFiGqvF7vtswqUqQ6l4ly
ty39BMSfeSRKptKnBaF4J0haC6Tz/wydrUzg/f6dvVcNhUSFsNbKffDYmV+Z
fzqd14/XeEdS89BF52+R3207uNEnM0zwPO4CFPpQ+59D+xkYDkWNs3/myT97
RPZLqyz1BS625jO0ojju7OBlF0UJwJI+p0s6ZYP6Y0+WlnLJsE/VABFDX226
wb1/NQhoaSOPMN5Bv8rVAq2BnBHDySHIkiwiSp862Ih0ZB1WoNLI3Vh/yB4q
uOD+ZR/t5AOIpz9ibtunCT7DktTA9257NfbjZEVOYnnp0bkSdebUcIzSOlH+
dCEn1qR47VMYpx/BW9hfMerADOF8FJOFPXN74WWwx+bYPawlxoSOfGm9lsST
8w7RZIZHfCPRWtqQEs7EZVH1Glt2R7OQV8rE/gWexSUJ7sp5M8nYaF4OQRI0
xpbnm0ZcDwJf51yQ9R6upFaYvEStoGRSpb7YMOrbb6BnYtYpBQ3VfbAU3bIa
23uxxcWQYhqbSxQc849reSd8eOiBt1++9szoOqLJMoYBd3YpO2D8vk3XeNo4
nGblanqCJzw40FOCRoO80N9LDsFRaBOvWyp9SrrBTgzW8on4fCjEIBggYQ+r
f9qAuzFZxlAH+GLmFAK2VSR2Ay7Eor4HapWDYkBSgLTngKrYD5LkG2fbINSA
NF0B+kiUEXrJE9XGs2p++CZtvoda6B+RoValxxjQdQC2MjIKaASnBKeiJlaa
ONKSp0r+q8BwZ+lRNf0Ru0awa+kxGhSoGQ34tkRQjXoGBHaA+G5NZDqAHgj2
koO9JQSr+/HHqFbuC2zVUdo4Y9xWvgInJhN/Zw2KE2mJyHdt19C6u709lWhI
fUl23sdSgXd0K1HyWIAycm9QMxDHXU7aHz1qFYsLLHxm0q1b74n9wGyNoTQp
7rzQe0oaRVyDBU6RR5/YxR7Nrxmlb/WLSBhTLSwng0a5iF4dfeMuo1sazIEm
YbE0WlNtLOzvhnh+9U+0Z7oiocwKVLkJpzPNCDPUelUdceUYwkIkduZY2r/2
UdgiIEsgMrsDm59ARz3L77KecSoV1LSnvZsl+66vHjZuRJWX96fwXmihmoRm
f57p8EN98qoet3476deFYg3uUUHOIfPwlRod8QUGIu1og9tp3S9Qtckttm/h
d+7ClMBFdIFsKe1faw3U3rW+3HTVjuwsLsZwg2MRqZzlnWBdm3lq3mTjJO5T
q77OKxLHle6FTLc+akOqGQMibS+l2iAq9S09bNuL2k1MBbkimctR0TW2pAXB
glVmpzSUj4avb7q7XmTxPblwmgu3JmiW8Bz9mjHWsKCi9favOWqCJHEr3wQh
NTeERfE97jzTzN1FI5ELgOoy1qSRRKwx1FGfFFEWprPj0qlpkPugP1D9oNma
d2mm7inv3qIEW7X7iP1MKZXoTKjAp8tiV8hhBFcjNEeJKaYeO4QRz9UAEdb3
A35jGp+p1IMViU+hP9PPzi/9iapcmf5UoyxwaIqR2Gajw+2OzK/gv/nUrdOL
ZtWXzWp4Vhobic2YiIPjTUnA/SWcBobWv0IonEx9eSlKcAYKxbYROpojlTz+
nXmRb5sMPL+AKbBh1ZkVy2GcP35Zq8V0KHnZ2trODtCa13ylvKKlwQKXadzI
BLdzYX4XXS63vN+zBk/yDiIJ57lotTOb4dw1uM1xwIwnUKRdmAAiJKUt/km5
ZesBS+s3EUkwc/SE7lFGUeUh6vTsVX7Du5zX6Yi8pcyTrP13EpVrXCvpm1cJ
vnT1HAF5z8/6sqXPNAhCtlLwA345KC2V1JrwIvTK+Z9L9DCX3JvkkOPI4nvZ
4TjzpviK+NS3ESeYrFc16fWIW/L7Zx3fQrRSCkjgj4pIoahe+o/EjZCqunY6
P7Nrkxi5j3u6epP/sm1cg+EYrcpOhJPjqk4KbZX0MGBkszOYfih2po3tIhKS
hDGOzGvtZGJrsq0iRTGA/eJ4RAAtLF5qFH6nbTswt41bFwJCG/D5bPOF9ZA6
VK99G58xFEZGf2uIwklR2enOpMol9tgaiCmq594mgU1AKxB4QHtUnOwgITWb
/kW4+ZUJ8nGgy131Sj8rsFj8AuCCX745QLOkq9nQEa5x6um1idRS/tUh5946
gLPxtP2TqtdLXPHQPK/lU0IbQq/LfwgdTzgFaGB1dmAcQleWzThhcw8RaEnr
0TxD/xcYg1p8Ds9FC/mPROvuIcbgdJ5nGWDA6akOzPUeg41bmOuYPhmOxoLJ
LkYDBCGGKpAgegdZnj7G9H04mfPImevWCWjxpWFOqfJAQUbTFm5BrC7vbcc6
ykdN5ANm1WU3DHgYEXP5VL/TLBaBcbrXX1rs9QlLJFBDQTvwvgeNuKYH7mYy
eIPEiWDnw5h3BI3EBCyYHTbCt1y3FtVp4QZ3DrFISVb+TJ0GXf8CgPE1cdDH
1bafGp4aOdH2jx3cPlr8A7dd9UyrW+8LZaHuN9fczmtoapix3KmAKOdC3fW8
rXoYA/nKYY1aqa0AvnPngFLeypK+D2QsSb9Qkgm2cuDgBjqTO29DgGh0eCX7
umvslYCFBLi5kH2QjlJkYYSS4+AZmRfmMhhLE4GmVvTKUiGPCWGznMJo2n/m
gXXRES9k9LW15xTDstGhpPVK5NWWD9tsD1UCnzXYRLRN4gjWH0/oevhuWt1I
vX/j6MTrouDGL80pY8CFlDPwti9yHgpUtkQQi8uSghVZk/eqB3cfpY5ukXc1
Q4UCy1maHjwhF+dDqZkz+ZBNUE5n5Yfm/Sbimyq9yY0LWx8GAYkppb4JljoL
mTSLSfX2ZjuKvXEKOIeRkGP43aNhQeUU6LKaY8x+kFihf9jsNcgb+2gySqCt
ar3l4d/SBWVp4/0FcFAoesNhmz5UMfxYzg1ffBZg5UXRlXBJYCwa1UXhxxTY
o2Qaa2cGfLr9a75h7ABq67FWT0d7ZpN+JUbA1KLqaaPuH9jXj2sXii76wQfi
yMHskAG/VRTrElPkGQmBXadFBPPLdvbpNtfBIuczZkZRT5qSQF3Kg1gsdGAE
eD4lfj2KWksrtYiTetsbgGl2p+ZeKRAoyJz2zLODmK8NkoXGnCO3eV9w5+8c
TKbk47IMUJHIgjhoOXTXvVX4NYtmkC+FOxEP/cUFjPb9P/yaYKAf0ExmDhmp
rFWAWiQ1SaT6mTadsBqv7KOxV+Ln53JJafwnxqF9sYfhmEg0JYl5tJaNYTCQ
nKPIzCVgPKE4WMli/wJnKyAwp3hUTZiP1nlWB7FY9YEFf1hTeosm9UWDNX29
YOWJQzsoV6gd7kiSGwHwNMbUp0urPDCYtbJBUwuW5/z0Zg1Uc10I+tdopAfn
ILviSu5lyarH7+UfDGiaqa1QQg4HEzn3Wc5NXjrpLuJerWz440fMJPJXIYQG
ekDef6mHxFjmdN4cgNBN2D4TyY4hOdIY8F/sI+9NmpK/T5qv16OFWxz49o/X
LLD2w+6NHPIyzfQq0ShFmrdwHyavjQoW9ea54TFjacYVzRPOnIUNoCACIl+Y
KtPUp9lLjpjZ4TBkM+hxO8hW+1RhrnplTXd/RreSp08U9LtCtYqf7/SsFY4H
6d7smKxsxxsUY9hfj9rWl5k4I+rgZPombMt6aABRoJ1z6UDWKaJBd7PQvxZd
V8Y2Sm2x0vXEM3nXa2dblsMms954BFEz5c/Z97TUaeutayQRomb7MgIW3ZbV
T8G/dferoylcwKjvbHqCqEJ0BE6+ktPpfK/oHkDh35kEYDbnYemYSBCJecPL
GikPc1m5ms6L+QCO2Ey0k0ph9CAugZTO5mqAuCq2ZnvJb4S0Bjc8k7WkvNQi
ZmOk8ZBM2NrRd4I80Q7xCZdl0RcSheeUgLlaBJIYQ0+MCCzQJddbIecMcl0U
wwaI84IieAfhFOXbS7HOvW6yzLR+zZIkDIvpIwuDPFGHl+Id7CM2m7rBldyo
8t4y1wkbeyV/3poTepj4SIwdCpZIECHWcPmIG6atL28UQJJdt6Ig5mNdjD5T
8l61GbolfFKWiYkQZ3W6azonZgImolL4noUSS90Cy2wxfyxeCEsTprr4sfMV
bFwNkRiamt46o1KrTyYayJQgpYgurWKC1wIR5q14X3qI4cSIkdJRHcJm/bc9
fSEoJjpyVwhHsRC89pfK3kSqUH+cf6UsMyQfY3s2pNUx8kNDSz509fGP2V2Y
ojgLI7PrkGaneKgiXSPDQBEy/0nnnFUEhtbOzGwfm3DKeHd5AA8rmU2ON9sS
PSeNnP/At3Y1bQkjIfMxHis7nZefHfJI0BqSaez6L5GvAIYnrk77HjwWC7s2
jTWNg+lO/lwCGPtYYCUn7GKNcQ8vzSWK4r166lS0Co01dzVlJXBaOJa17lR3
/bQ/lvkT7FUCRr2LeIoNlG+m4PU0gL08/gqhrSzOGZI3pnxEZ02FTc/YIY0y
i+R5daddNvf51pQv3uiJjvDe8cbfENMVPHwl5dYoHrnG212CY/OGhGxzQQgD
KhWS+c0gABRAkkfEtOVKww3tmWjko4Mfdf4pXsRyAEixfDo/u7vwnYf3Ft/2
gkQX/uuab4N1s9eqYhWRjUd+i5wU3+kz+RA+mSfy4XixZAd2GH0sG885qYC7
vlGqlmrKi+mVI9c4U9vpwPBGPrhrDBi9Plp4dlfFRz1KQWm1DItj89QS+pdY
eEBFygKyB7in/p4QRg9YhKfnCnw0QzapAXxuwh79J0PVcLKkn6x+s11iiDWP
RVtSRS/ebw/gklHJKQRkYHt0NvYVUl7Bj7Yd2WZ8jb/Xucr3R3RvaBroXxjF
Em/VGFyLQllP7fLrEoPSvNqtLaHcLEAdKIYLam0xAVbuNqOjRyCLNyxK4HoY
/GfKXQVVs3NYGdDNQJs40GJn9m8WBibLMTHIv4txnN+zGpiOXDm6m8SS5oZP
S1WIlPD/EaFTdeVMa8V1kofIw84OqWScK3Y0I5XcYsnZaf8BOu2tCZ/m0S6j
UqSj4r4PtA/yFAyonpuIU8LL5YhPQBEl2wpD2h5w8rCOFgJda7fms/YcJ3zl
MN4vROupjL7PMh4mBqLfOysZm/2J9pVHJnris6cmF/pw9y3KicwoWoqTm6ww
5J43ppT1IaENZyW0zIoa3q/723Hz5G4CoOImkSRbKBbUD/N3LigG9uOVGWeH
5qzLA8DL2IBz3zHyEqaFb3Cn1Qx4q8vhAJrXqDLBffoe9PKFJ6U9EmjjFK09
XpGUWCJKbwEKKvH6oWTS9LTrt2jfdWWBeekBPCUDDEvIY3xuZrV5YnEAymdm
4wWAebY5yE0lEq5nYxs2xg93zuSgtm52U/No20bx2bS4ifqQXDdsOy0RIkzF
+ImhxiVqnriFpNfknqq9R5SXMq2FBEI3b36DbbMRhI5/j+xNm1d5mYT5IJVk
QjtMrXW2mLisv+t/kNu/aDdVm8rHPcfv3XeQoBUR6mBkxGTjwotzcTUpxxvR
/ARO68jXgcgoCGA+9DCdjJKeXqkpuV4PD5dr4v/taHwiyQqqsQqdyDTyBcd4
8L9i+Tid2I7zq5M4CpSScgOAERyArTqxHv19clXWN1+7c9BTP+wD1Cw3R9nB
e6Hn05BCajlsDl+U2bAPtzGLVK8O7PTI2g7rkEaKAhAEAp3WK+peDiS/k3HL
owg5P4bfiPpTIcgjRCl85VZRKXouUOsHv903IgI1Zg6RyEnc+QmDd9C0mBHq
SiiBFQZf4VwpkoJ1YAR9v2+lCpny2x3vUgDPcr9fkrepnAj761G3DUP+bFct
hEl1deu0UjXTDeBhPk0oxgNOtZGUyRzSRsJ15ZJkL+7afNW2JjSGOWeyfw97
gwTIosuTpPUV3LFCUEnava1qWBeZwzS8EN9e3vmzOzOc2y1lvLeteqFiIn4r
LOQAXqL68heHFh9y/tGZ6KiSxRh3fvA2nBrY6/wAp8wkWq/lb0hzJ+uNJPOv
u+Q4ALNsc1BAn1lZh1ldVIwdibF+8GsqDrvHHBIdzXfLCjA+w3eZp1akcg2S
oWdIy2Glcw5qO8HMxcKEjZsKO8s+kN9Dnz7eKhOuIE96Ol9+B1GHRbVjGWam
mwkIr6FnW8F16JMRGQgO4DKKBGljOodN/Xq3TX7doOgYEzK8JEC2ZWHzqiZJ
cgW2tD3yCVLPMvF7OPE7X1PDRYrEHxvltsbpgJ1i1szBaMYxcA+vxluNQXUb
1nKzuOluu811DWqfa3TRCZ1tQUFJFfowAcdfevnNplpnr7Dxj+geExfQ4DYD
YV/9gMDoSGWQYOug+U/rLfLYLrn7JUvCNjDtO6OgZpYwWyXoCzPzpTjypTM0
T9nNRah/dF+VB8fCZtf8DV0msfXst5WfEPnmYvu29PUBtJNtgDNerD4R9mmP
rLRnkmWX9qePCuWe/GxcAhu5WRPrw1Q/iyn6r5okLyF2z6qI+XXoAwDsLM/p
pIDC7ldh3vPmpetAP9J727l8zZu5r9hrjgu+hlFv/3ITE2swgW16zHf0/IKH
kt8cE0uXs2bwrgXHo2VHqH4k2cdU7woLSvXE2QA39m2QuoTsF7IN0u6VZ3o9
RPUwJ/oPue2lteSOPx+262njdv4J2XFzNxViDOAOI9pMQ0HrkZi8K5xinXNF
yrefauNu/8iGYhGXXSIlGmwuvjRIIFFSRArtUWLHMdHJAbCMMTGWrCjHpP0E
M8kl5wi8wmnTK358/GDN2C4z1aDeVbBGU4R55daHhngSA85GQ0yAXNHOyPkP
3xC/NLfdnu90aY5jlDM4I7NxZNrvWkQhaq7mEpsA6E6Dcm/qRAZrzFqKK+UX
onckU8pf9O+D8P1iXFvmSkq71JypXkVN+0bGb3OELPPrPftuov0CLztNPUu5
VN3JEj5ZheK/xWekNafkrXvexNrGw+2c2OuQinLISfxDmyPa8hwZn4DxbOgT
d7mSp7kILRddehFmaauRf7mW/h2awQbLo8LREvqfd4m/jHRHi3xXuz6rsRGm
gv2L9i/QOoNrt9wa2XPusalOR1fW0naKxRTjqyBdHtbIUPvmd9fWBloZql9r
0mbJ0d/ww9E1DaxuG9dyyOzMR+YNRBcO81+rNeUuDTQ6HzVcZhAsEGfbRouT
bLs4813sN0l6YV4jXxfx6yzapl8QxWioBXexeuiL4XFHbRTPbbLh77j8wzqS
6QNUquDrt9b85a4FdtJtjZmbKpfZ/MYowySP7wNZ0kWospZvqEXb45beszGv
XShv24/WtVYyZi8sAlpBk8SEGVo1KCCxbGMKZDH9RXoyvsOjtr+KbSa3tZj5
5ZB+yH7sA57G6KusodaxdKv6v04Ns1nybD5qd9nVAHwwYw/cGxF7cNUk7wnm
nniQiI96lR6DC1/5VJyGCu+j98UVL0otQ+vuUzg3Ur3lTnLCLNJ3EOfBlYrN
K9qFoyUZ94Xo5uuRZBXbdAcnawJQFtvODvBXmm9gdTXZ6bLqddfUUsUxrs08
4fUCicDO1oUnfDos0EVSobcJlrxrmaykO6OA5ovcMCjPT/iQ1WA5KEOiVrIB
4YwTqBPrp6lbCpppSj94KzOAvD8v1QSOzM/MF7p5b7k4UmiqQUDlRm9h4eH8
FmoQ79hNhuWVQub1YsFXnffB5ws5jbEVHNplgeULxVfeex8Dpi/BbHb69fSa
fyZCke+/HpQu4Bdg+oc/CsazTbUbPvmigmn6MAfyNj9Zec7reOwCcrSFHAuk
3fgjrlvonPU8obAxUxcKll5b/s6EEtzZXM3WYw1KSkQh3BuhfRFN30s8Ov0q
uC4lcyshXpF12Ll0V+gHDNwZ/FSuQ7R4rcUsq6soBSk46EkfhcUdlNGMC9ed
d6iv/m8tGPTY2BNvY8q7oRceyUDNvhJoR7YXNKSkqyeF9RMoJrW/5vdKL9ib
/1UQUeaRF3mDcGxjForYyP4jHXbq+IOdcRo38HvCopSA25heHSkatS1n0f+Y
Uc6/4CYJydTZlwLbdLFVrYp6ornUC7Lv9/b97kSY3OcfQqIVycPFRqqzUOw0
z4j0lEURbi8H1KlkDEiCtCnSUFLLsmTrJeX7cCqXmjKkaQc0a+YIG9XPWJeP
ioZMYqyTWPRoUaDcxk/7r3RqfPdUocUi5DrU6Ix6/yD5n00TslnFy2WyAKyu
hRIMcpB3s49JxY+I2r8x+NEmQCNXJDSpHiLiHaXvoziIboS1uIf3GltvXdCj
JhPMqmWbQtyOGVoZzbe4JvngTxf40BPpp1MygHHO/z+wo1P8SkJ4xuyWuyPy
b/5hN8fsZfQl7vCSlPR4mH3yv73Cy5Oa48CeQEIR60GEhH5oh1jTISsFczPW
P9JoptdRxIlpTLxcr1JJD+hAP5P/xEkYQsbcdzMw11ZPPkCbEDd6uacBtVfW
C10G6lOaV7wrCNd5LuC2FDAqZg6HjdHXrUkflN6vf+BJBDTm44ORop0AzhPp
PDsCwvZmn9/Q401tkSPEyfRiceER4RsgurUGDtQMBXtl8xucTRBOm/2ePRsi
P1hUn0S5xrfXjFGHDzULy7OexPTLByy39Ww+nv8pRG0N3To1SNCtNPar49Dy
zTm09SzZBsLOIAfNByrfxRNXqHjp++GE9l16nLe5NqsrzvSalmVsZxD0c0Go
4fnj5ViHNJH7VQMvO+aqLyBvX/jqQh9LKotOEABnnRdR8ybqeSF2ImEI2tEQ
C+sdDKIXQVJ9e9VB4ewKkwGVKluPVct+bsndFkCC3p7/aZlWfXsCY+64gfda
hEZRnxax06iIbtEArd4iV8tumr0m86LHh4VVYZwDE8KsqnmjTcQOKSbNCetW
ijDPOVMyMtEvZVMoiT0w6qO1Ecw9/z9ZdpAOiU5QYFIss1Zu7TFy13PMUY0W
yk3uQz/4XCCEfWfx5zFchvaltSkJUbQx89S4M/hvjD4KGaqGbsWkzefyTlAM
LuhFb6TW8+fvc1lmP3d+IrPk8LMKqqcwUFxf/ag0FICXEPw33Cgko3CpmvLw
m/pZ00KAjB91wrsEREACeOhFEIF5BQKprklqxGqUpQeQ5QUVfd+FpOLttXHr
MKB1WktQ+aZObkH73LiSNqNkrE7Exg42pCArFIBmNatDw+kv4IqRe7w/coe2
ruJ9y2oFtzW/VwCOhSLerrPSK6fMd2ezXurjZkRJoJp2saopYRtnBEFoDxxI
WTG7/wcx/53n1dLvg/woaNHy8sKkJ2XINSACSdhru1jHeWxFP21mnMA6cRMS
WQUVZaUAu/zYhA6a72b33zyJJTo3admOnr7RebkUbVNlDuTWywbK8AOUB1A4
dSBsuNcpQrvob8l5YR6kowyLmON1opQHP3EzRkHXiHGU/F/0TMk/GIOqb6Xh
lpzIHu9lniUL5R9I58MN3A1nHcEUuMwvV6z6/aUNP7fdH2IjjBeC5cI84EK0
JZVBjXjMivuXog6qUH+w3hnXyrv08URVsuxr6KAEe+J3zEDzd5/aswSmfn7R
1vV4N1gsjDrWWaGKFIg9eXoYol/XQJAadzoqevrGA7nxzYkoF6PJegn50Byk
sIr+4wYEzmu2S3ChOoQovJpCuldOEXER3zUzKMlOYeQp/nnbEa9nHzMtkjYq
O+O6vc3nWwrn8crIuErfwwterT+Lk56ThEmtic8avMvpnHMtrfe34nThSCdW
6GLOZfecqf7uHzraJHaQ0p4ej+obxv2BGVZ4p6d+4zgaCf+G46C1rMlLrJKL
jQq0gA7qFxrRD0q06IBqZu+joqJLbYQPPVcEiRedL2TXIoIDjWmo7Brsw3Gk
G/ooWQgXxLYRJmG8G2e3Lob+LGrmpLCbgQoyFPHlK7BWNANGLGQ6OjXocXwO
ePCVi86EOSfNFU2FyayCaB6b63SVxkr6UKiohqixMe75tPMlw1VdmY/fNZ8B
tOTV5XSK3e3BSO2cgArJLxVbPODAPbkT15rnEz7j5hyMPLV0A+yIv7zFPr56
z8y7p+RFNLKFgxy3Lq8yp44gcKahN1mU04gcL97AeI+Q6AVLBDeWZxtWKNEM
XoRFOhjOt0M1dU9DycowR4rnnsD0eVA/aHMmcLTXBuiJzP9uGj4V29PCbiAR
Hd3DuHksIoIR7WUJYEnoNY6VJcTJg84a+/sU+Rcxnp1sNmSGPfFU2SOtIBMT
nANBhx1g3zddqyXj+YlneDvmHtoNDwkAg45sqGUIIueo1rmr28oKjO+lJ6sx
t78bxWerM9w70BYbe2T5UCQXxBVVB3LyVWTrZXWAXjjHLwh2+FigneZ7nGks
achZe4uXUmSL3uRZxwKA/3TFN8sS2oBjPqoWNWt2++/rYpQ/qu4CeWsOqy2t
CHXAhbbc6zKgpLLrnFsCCTYqxE/DTsD1C0nYHeh2F902AU9vdg/MZTHDxeRs
COg+32RcmhM1h7yWZtYd3CtrNhD8M3KAA+3xHTNeTfN9riLEA+W/lqEqqhKJ
QyFcFo035ZNhGQZMPwU1/ESh4ihItVINgWvJuwXK07u+qWBsJEHoe88WANZG
7fRPSf064Afc1nxip2iu+HlhKszUbFsjfeDoqGk/kLpPF0KmOVWw836ap/l4
wsFdrVvCm1YI/e0F3Fm7hDx3MIC9cxHRctvMrF6hdt4OasQ9CMLxo6wLO9Ax
cYmdSkg/cHIhMstRwoq5MyRjNZSVdzgW6iHR6O/xYFDRhYYkgRBMXZ43HABd
BFqx/n1v4FMY26pW/LHkUmJWu2gAMxX+MjbLFgLjvI0NprReCKBKAVpbky0L
Y2urf+TBEGoD8iBCwZIJbRDW0SY5KoMy0GYU1vnQ9l5+GlvybiJiwjnsxp1U
uUg7VONymLbE8pf/s6L0vW4HSa2saw0kvkYCZRmwVSL4ldCJPghQ2+ozSQNY
BoPmaoCVgBIuR7xTyGQTLDotmd+YYPnRc66Ydj8hQKyGWzB5cIyoc1K6dB77
HB6I5rfAndF5EQZVWW9S7dT/00ldrBIjDas7lECsgwROOz+LANnbkKUg6NcH
Eq2G64qdJ/z3IAeURYj7BIrQ7WFDZaeql7w3wFYrv112ktBDhtaWR4UCscwD
JuyCAXNUoBm4KvmsHyN+BFZ5tvuelWB5JpSlv45S3ekZyYVkR7cCieE7vMiU
CKh+hy2NgJXSapGATvVFKERH/31dZMDpzdbI1imSUDJTr5hPatZn+5jY/GCR
Oltzni/qWfYOYs+aZVttYasrKQk7UI0GHoVhmvWoujmPBnFiA4nr3oQniNV5
VHf9FTNwbMaBgN4QcnEkzDSXKyz73+pJHLnABtWl+P96aM599G8gXT+9+s+z
/NpCyazn4pQVVrkzez3zgA/iPZfIRhqhKcAJEUhf6zAnAJx2gKVE1i9s6+JQ
M6AVgbJ3i2x6F/k7xHbf8yUnbZnXIAMICj2nDuIaF5/vHUEW0Hn0SnE4ABz5
2hCmEuDMkS8IlEhz7hWrbSown7XjOmt+eGiBya1mTZtglSYofbvXK0WSfEqE
tbmIZQPxdCg/I2rdnrvC7GkTVPdm0lbib8huMqfDC1H7R029L9OKjj8vvdNK
m8kncvy0IIIwOeameAxFF6qGkkZh0R0CSk+Wn7+YNkf37BoamP7ArLiMIAh9
GUrHG3TrsMi3JIeWmhR0+0FzoLsAV4+Xs01rozGAq06DiEZcs3NgnctwsDa5
67Rbni/CyHprRfMbpUk6fxvDvtOZhUkCybDnnMJd5sntXLENy9TAJu5rqMTz
oVhNzopyXL/5vSWPeFPxeMRmikEdOR+e2Zc5A3YiEX/DfXkA7x30NkgsKzoI
Av5JciLfDWWKJr5G7v9ThH3ZXIvESYwYTjhK+ILGlLOkfH/G2yjmGFAC2LBv
JDLe/1mr+AaHO135m5VAVdLgQbad8JsJPBGH7yQLy8J7/20lsjT18INYDDpm
HWAyIW6azzYVjXFyQX6rZl9yzMCGtq9T7I6fClQa9C1HAoVmFZ3QNth8PqoY
AP8QCPTDrBZ/Hrx+RtDJznO+9G/6n7WMA66oXNFmR1f8n8hYlk3qDnTb80/4
yaVomg92j6N/ISit6av8TzrGwv6tffZ+OEEaNdBU4zxi1O7ibwsgHafnzXFT
sNEHHMFCdq+YgZ5ZTc8e0VEpNilf/WhDLH141cOikEyUtfX0sbLJeGLXlKZ9
zdDVLmA0LZam0xBx1jxH97K+AWPDtmOnFLqQ/SPEpQl7lMQn3CBN7TBex/pq
NA/rbSveduvZbYg2olVqlCC/g+7lvOQB6+FFLxpG3WQwotKrRYC0GfMw1mKu
MESQgdzjC1QiPGTu8HLTq7RoRu+KV+yAKEv80rp4mfOiaxg9oskmStbID6+k
sIDxRJD/CDNj2Ck7/PsSvXrzV30kYJevZCvHAPoIraDEEJ9zlDRzm7lQIS1J
iguPq4+3i2MQNIxIx6jw4ZVDyy4pzoC7D5KmteTgjetQcbWiadiwsPBxQYtH
5Y5VENAJXRKk/BelhPdsGhu14AT++/Pph1tj3zVH2pLIq6SoAkIXxE1tVu8F
LeKeEyZDjuyofb2QTFrNbWPMHwqVmlg0XezDThWj83TEjnTxYSdbhg7D5b4k
gLWxSHPqDn3qiGgn+xOtLDX2V9YedrKutVmnbd2p/L18Behpw5mOBCq4Ukdt
5u96Q/ljTPDyH3zeNmDnqJU1xNexz5Nhh0Ijg//1I8l9F3vUWAiLsjkgue4l
sVrr7766Wgn6OyUiq7W/EXd4oiJykZmhaiFNLgrQvT3DKQd8tTRT8YjWvmEs
6o41wQNc4UCcafu/e2mEYBXnSdDdxTzVIkohgzTB7itQ8T7fACEnufQFI2I3
w1qvY3Z6xei/w0sklpZ+8mEPOzG1PC98dD3S97K3vL/TUX35nAxSBIhfEBCV
lKLKekGYhUVnZyUoBQMqhElM3iV6x5TE3Bb1peK5Zx/5Ffq5jdFD3dl2sP+w
meEoQpdhz6xIUjuGfxPt5cIbTw15AWt499ZIP3ePAI6Ee5XJjFvDPll/hwXY
dSIGFUOqykFFx/mZfRiridM5fmn4hAfRMRUZNN+LrOlmURewAHgBZmisqZT+
c71T2js7AP4sIqD2D03vr/Xu7secC9JT1YjLK1BdRYGx+XtMGZkAluytwclb
a4yyr7HTKwnBx49oq69g2XbuAePHhLL+K45JWolefVIixwDin63mFmIgOmFA
TU2qT9leFQR3PHNN2N708PfaHE/bpHDXgim6U1KTjbPOe2g4Rpx1qPqOM3Zu
JnHqwZMMhNtceJ+3Yf32/xj/h0vu/RIGdMmeXS8M839Fe1HzjweHRHhG35uU
Elymt30w2BXVRk5kyR69zxhhxtAd6d0eLH8Rzpcxol9LJQe2SILGct5ui/Nk
ue4Hb070rLobAZmnq32AWj8KISNZIFte1P/jsR/oWnaMowTFKaRplZXK+1iE
n7wE29hpbg5e4NalPY6RbSo+WszmUF0tiQRnMwOlZ7BDiGorJoZpeVwbTnx8
xDOvshlJpireSjq0a120kyl2RsOfIr+SoADtixJUgyZKcbmapc4OoQL1FjQK
WDwxzzSUAm2BXA1669c878xm7ivUHuCwAIpA6axivJ9q5aGOyk0oG0yq73PT
M/4YLQ/KMCSqZpAb+Sw0baBf/9yV6O9zwwIIqzjCPCE9ufFWsnPSBe6kdVgC
/S6PkCdVVHx1FhUP8CbNy/FMVS8XuhlnJhRwANYK0xKuVVZM8dQb4nRGtRyt
9JT60dNDO+jCabt4CpljjJBS4OhZ3UvTjL+NQQdYTy6Ijbv0TUlPBnLWPVzu
rk3VN9aSan9w1Nii5w0L5O2aVepISkxhIwSZnM081r5wHbVR18zRdIqj9zmB
KG3bgTsY9i1abL5YNAalH0OXlQ3SMdu7dCVmiKsGWXsLAlz60qcu0Mj+xLnL
/CX1NT/co/mSHicp0URy1qu1mSb1yr0iqocC1/NNovLF5WUFw15A2Aa0JJjd
KpmdxHs/ktQo0H+kKHyNdKaHAh4tTD+3rTC6quxW/apJv4ImBC5ZgskLt6b9
oqgNBVBB2Sns/AlOr6E1xdXEb5hN7w9/fA2h8uwv8fsaJN879ktHnYLA5p2v
WvU+2IP3FtRD64ND9WwWMbK6VXKSjTDHq6ule5F5wczOHm+x1Rr0e7N9IG3W
XsZLs72DGJ2JBhx1lvMDJWqPvd12rm6MvMkO5EjdXfP7kGfbQDYiMWN3w2i6
PHi3dmzCz0fcz8AqDw5iK/noFA8vhyISS7kPO5GTpVcMD/6R2yJqdFB0FtV1
zl09sWPYZ40SitiEhMKKKlkKit2qpuoE+erv5MGSbuHNDDPY80vowOqVXTbP
Nl13rgYG0dCXxTLz24HwZPAvewVbQmToPNHGxP4KIS3cklZxaZfuPYCBxfTq
Y97PxIE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI3FgNNHBauBLYE/7cqQK/sCnsuOGE3m/UrPI3b0iuQAP9nKxTt3CGf3vShuGoGspXCwZpUx+YBLWt8BbwyzvYhLYw3sk0RAkkeKApT1ocQAA+gWH6uIF41m6htv2aVGUw40hHlXg8wnRaRF2hh+juJ1mEWiHPBDGIjWH/dc3HyfceItdJ/frhYvCfY03OFpYASSddp05EeDfoeSOHWjlgWugbi0H6e8FW9kl5M4WIRhVcAl7PZM/xqTFNuVRz1ImSxjggI5IXsOlfLr26jEHuo1sbrGrM/KmlY13IcGTJ/p0qjHRjcFq4Brt79Ap39Nts31d5GkgLSJQaz4NMREUZ9d5FGt2stMXR4cdx7hH1BNDjHNIoDKTUR4Pk0cnOAbQ3dNbVQJS3Efbjp7PPTPZFfxMCtEarV/nvbb9F6UcO3WcuMzkULsFXcHH7rBdXjuMMZpjslVMtwNI+lbBkd2/2mSzwbye2ECiKFtFeUz3voN61dic3CBU7vEzWZzNV7fr8kcomg7B9oEJPCLmz1qxBHukQdpMZsXKM5XoVjEVeYAPN8VxiEGzBI3/xngzEhOLR4YBt1+fSFpgvQ7p5mkgydpo9kmI0usgDPrRP0LT71sBTCNlRAf8QGMtrrA6ComhetFld6iCQHeOkdoS1mZK1/PFRTNVPoxu+LFfVWnbSrWABdF8DExIxy5ueHBriZXcABjIK6vIuI+XQrKu5UlhJ5preeDgNuf6aChTgxfD8Wv3UdbHmdEYer0czYMERTw23pDwsvMt/k8rxKHsSaZjrVv"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Suhoh8D7GGQpOjd+UbvN+PLehtn9q40OKJaV9A9PWTdUZcxAlTrvNFAHUNnu
p7OjZWiCkU96Ig6p3ykMTrnDI8/p46Cz8G+ZCD3/lVkb8N1+reNakAUuzV9v
XAkC/SQHa8pQzxkc5ZRaWEMTF+oWX7yGcPcpJxOOgsG0XDRHB7uGBbjLov/f
hr3sGWAc+A90+p0xYCDqcYplnTBziXWZS86/eUxWGEZPqOov70e/9uKZaFya
bfhSX2emVvSfiEcUpiXOzd5TJIozKfoZQriX7jpEtH9oq3z39ybdJ6Ys1iL8
T5QxF+amQGurWnm2hzmbF299hpp3s7U+q8R5JV+6Iw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bY0yNYGP9fUIX1RaZ+0kLiF4SKptk6vohsWmUBKgprQq8Ip24A5zAXbuEY7Z
9C0SMF73NX6hrYhxpdM6DkizZue16nnq5yS8kQWcTRP1U07wxFyGK8t05MWp
qJxtMMfskdTuPq5E0oOI91gCvNaqXzXqys90owJ1bgRee+2gXDSsMj68wd1f
88kXb7qSa9IvJWDhIeUlAx9dYbkh5UMZSj5BzHb0oijpTAgW3RNLCxzDlaIc
/Ylo8n2ZxvhoSrJfPB1n4mZX5hAXf+0Q3Hn1ZWhhNvgH51Iq8ip8o4tO0pqf
XoFJNSFsc8aYd2qVST8Ny5wOAgD2PvvvjHSzWHwVpA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AcDwPMsM1cj7bd/QdsppgW6seiHUcBccUsXx3WuUEVHpS1PVMznp5ukisEYu
dtM5HGe6KJCnl3UL6EW1Rn1RxA36wvOVegIh8dASL1LzkBfTEhQyOVgmRKQr
iCuRvARDVxJ2ppDKAWeplYxjigXW1MVrkWv6x9JKfwXKZDpIHHSwVKO4jKtw
inMcRj1dPCGI4h4l48FGWJrOikuBxV+tWTHo5V9JjnB5YEQAfFKD49GTF4wc
Avuu71+OQ87krF3V+hLgn+lKTlnigOzOlXZclCTlm2JxYQ8Ydg8HrkzQL6Qb
JRmkwMqHXy1Mhvd0jJ0RT+hJ1pF4g64sPFdxB6GzgQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g7mqQILS6T+U7VPc4Y3r0l2mQ2NHzQzF/ysxj0aupALqW07FSgwIGfgUdDof
eUvbcb0vggmrSvlExyBnVv681Pvkoa4IfwYH9Ooqj694x64UHDecLDlZzNO3
i0QtNbQZ008xyuoGNAbDeCZ71SFprfx5xrEvaMWYQmOTqCe52DTPrV4mPkz/
9l7PU2x219bl1Q9FoQUW0WzLWMFdw66ySINQnf/Tj2UJRWOqt/RuHcoHFc5V
2vsSbmfBgcB3kGcsQs4dDSx0magicapnAdEqtvMJp9yPheVyyZWaIl6QqjcO
JI20FuiloRUPDbRVpa61Hd/0DmhEoYImc5C1N0JtKw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DCCD7JCaaKVwI0kXUS2X50GRvLZMs+SQl+RFlen+DVwUWPah0XCsczyfqzCW
EN+87gvgjbZgLbKnm6zhV7VTXRZYyksidodSeYv/uDBtWpPXdm4yNJOiILBF
EHjfTqDKorkKhrepnMjM0yc1dlPMOcG6UIwTI5F4mqGr1achzlQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Q89sYDfr9iPHuVvgFg+EGGz9WZI+zsGUhKufxgUum6Ps8KYCkswA+R/94PQV
VaWwskKqJNU4RGHxUqEmZplaY7LIMwym26CiE6VIilCn89TPK2onx+spwdJw
NDY0UaqLZ1beOlMoEpbF+J5Mid9cp0WUoYrP6FpfarkWKLCyjyjhbyVo9c4+
5Q50foXnb4NJQTSGhPjAg4+J0j299VZfxKxsn8xNiqleZUhYSNpqxg6ERwnz
vuYbpnr4QdJzjsFyNdiFTsvkgDx++Bm6KRnkSvr/1zoLGeIcy0rk6aBcBoqI
bgd8xdGj5eLwU+teYa3m3rBcKcGLor1hBAQcVEqBm76uYeQqISbGp07SI8O0
45hxGS/OOKI1nZc4Y9RjVb2pEVUmx7/DvVi038YfAdGp5zjg9oJ2wkIU+EKz
NH779zmXltMuZYYF1RawK7tDMN1hnPloSdvQnnFLfsnuwtVTPYNF00O5Ja/h
Mi8iMiEtSkaXrn7Yr+K3hGAp1A99uqgT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U2f/9mPp+UOoMIQayuq88wX6hPkE5elE6+1aysPr82K5dmHzgrVzqrUbqZTz
V8conb64ouhVpu58VUutgr9CeI97C1Ivr4wx5LL2X7JjRujco8sAU1yhdI7k
U++xatNjnqrb6zdhsTpPSu8vZ9p72Phjpxp6ReX8neKa8vovxRQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qpTJ6mQPhfj2rrbEqmhP3/nfdFUXvRjwE1WONXeaKtikLIZ7/GtX6Met0E1X
55A4H3pRjTQd0L033zMIdNwNpx1VlZJakIbFJizEsmExdm6uVY4Yih5f/wTp
0r0nTrd5TnMMl2vI0FVB+yvzgfo+m3uDmYKX+4gPobObclUUxyc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10512)
`pragma protect data_block
/m5E+jIwenQqtfTk8xlTrkYeM2l+SLM3AII+apsb2qibZYh9zhFIa1gydwDM
ThDqC6BfdlswMMzM579YikJGlXiZfJyGanYBHUq7dw/zlsEQZO4BL9y1WeE4
zH33n059YKpXRKMHV6XKeJvdSHultpVuBTO7rNyR43Y/EoWX36CnNB7aqKH0
EM1Lgmtq5jxca5+iTXMtK5s0jQ99BQQTfihxFZxI5tpWyVP8STFD5RQkYhI0
WSifBGW1m+1bNIqENMNpjVLONVgflzYJvOkLkpLQ+z73OHBPN/27lpfO/gz0
QP7irD+sdOYMHmRygLIEp+vKUBb0fZsUPXqamHaaJ0NFlDAcpZO2khh962Zi
Ya0etmdbVU83d7EPzJmuu8FEdEV/AY9ZVmhcGM3RqSMb1TDvBZOJozzQUswb
jUX7WGiUUkObudKyJnSOfDqfJG5g0BWPr53R8LIiL1Kk8LCf2yn00F1dkxBw
sQA1myEtJEVmynCgwCBdilyGKzFfwOZCjOx24vvxda+clsdi8VUXzje6+l1R
yufCizo2HL0tKjA038P5LRxiDmLpggwBE54hcoHUlngErU14YtuZ30iv//Jo
w4kOBtuyuSpYmfzanNrmuqpT2gxHsyJKvOO97HgDSLOcki+sgAyUHIlbI8W2
2Repcrte6bb0zreKusKuSA3so3BLZAa8iubcdEhmrElbgsVxquA0AlsnOXXV
UQ40A6z/qJGW18WOO9UiRPlcwYL3z1iFTRrDUBFvUq38c3yRMwYF93pFVSvq
NXWM0kUn2Os2hlam6VJy8CLIqsCa+mGtCwp8P8KWD4aQaXecklm3ntg96e36
3BGCCouuWjW4ekG0KuCU7Ifr4ghg1F0pBMS1RyBFt6NE3p3YJJMkPny5Xrje
2P4qkof9NY7Uj+Zi+4b+Tdi9y0xASZVwsufV6ydrAvEPP0BczTXRNHq5kW5/
B4oT8gJ35jjHBhn5fRZ7xWqbDOCrDkvqCMZMWAhHTDlx4V/K9dDlDRSt4sZh
LkSoz/Q4JodiZNNMlToMP4t9mZs8VWL/RDw/Jih9kFKTIQ/OrNlFkBNvfTuV
05xCiwC8YAUeK3nEUxqIR0swFwH6VzsBExkDwL26+imp+Cwbx5FFayk94SGm
0Ab8U4ZlvHdYfm8JjZlFAvMRlp60WpcYkltNheiQof/yD1a3tHNyE1d21JR0
2G5HpZTaIkwNtprwj3ug/DjreJefDgq84cShCVUWRHa9eWS1ex0hQGs/rE3Z
jnPRXQ6SePrj4/98i1Ybv5/6G8itEoVc1R+RlvRZYAnFFjFIAuSmUUv3LodM
+B29F6lukOu1Sq3v0Z2GjjPs4OZxADZ8OjmkLazZ95N9AwwKv5j419NZ+x4a
p0RxMLlvFdckRw94OpUuEHJ+63pHlMRWq9gVXz36ji0/5YxbcLe4/Lqx/Dwb
J26TD+ue4FX/Kw+1qQ3Zi3jZQeWnIEdDdYRYXn7gmUgm7yfFwUpr1B3P/I3L
UyT62Ps6Y907U+FLCWLIrtb0i5kxtymmBKwEgKiyo948p26SPBSlTf6r3OOl
ZunqbmDQydL+GQZNqIqv4cvRS8HUk3p+pW6DfQ2ysLWWVxp+Rx3hiduSGmTk
i8pE4Eps8WOh3GzQjbeZQAlYu95ftrh+pvZpYiRmjCtHR5Usa668BsKL7pAR
nc/Bm58QS1+31I4DlEEy6RGxn0b48zpeHx2FhLHkouqJuGUnjawXKhnZjFOU
xUGqPVC1cH4VHZ2M5+bL0SU6RiUx8oj9zP3/zfpZf4FTJnaGrsNaLlzSI07r
jm4cnUttx42qOLgGPcRWmL8sKpVVrUpJOsj8GYOobQHlnZRfwCQl4KJgA5DI
Qwg7Ii0Ft82d8V/lIZrDYpPIOChfaYhKG7fMu8niDkWuJ+QkAr5Z/0ptX7Wb
WHBB4vCIrEreRs+kP+VOtTMPvSrVbMJjBVt14coeMauhflSClol08Q4Mc4R7
5DRglHkv2sWCwDumQktHzS8x0Yjd3wA/2SOi5iOpXSi14m3Iw4ynsTmx7HE+
OyHJ/b7nkQ2ieyyR+IApFshFFYAyPXiT74MvVVJ2/Le464VSkZ2nChkU+F/O
BGNvKA+Gyzm44ImtepM9mec31HlRTgrMdFaXDyGaTh43mPDKA+ECKzClHrcM
S/mudrHZ/w6LCVTIHepf5Cudg0nMkjY6YPUKYdnM2OTJQHTgGOhRkarvHfAF
uzMfzz3/qR97RetuCLHDwawRD6H+kmKa8gZ0J2gRcOkaX4BDvijILQnjuQpj
3zU6i2FVmUDG3OFO08Wj/T4n5V+xfdKboj3wX6O/2GXvteY2brNGqkMJAXpD
PkNIef9Iu44bnQtm0R+nDCbHzHvna1sgjPboB16FO6hzPa5Ntux95muSSCtQ
ETkrJyx5a0y1U+vfq/pBehEIskiVgcaJrrzo9WOzn52wmkva8s1zJK2qMwmg
cjWP3PEVbv/aj963b2aQjq5JEzxDP0VhZg2L2LjsU+bAN4ve3WlxWSmLZOsH
Dda0CEa508w1sOrqlj38OS4I+G7hQV+jwyIicrJD9X/Y/sc2ZhsiJ3ZF2Deb
XN1EsEaT7XTaeJ3v2dONM3WWzjbHgpixAcNq0AFSixDnI/PMiKegXBlI4z57
5bhSYIMj8LGkSrohGVpCQUWFZZbaicczy0viu+wR5ef0yGgOi4xDGu4i6q5o
Hd3qrU6JalCxVTQvckwIo+q4cTv0aNd9zjbh3lveJ+cBfcHdw6tzRZkANGT+
vICA+6u0PqO4p9gN2WQv9Vv40j/5UaomjXRzcmbfhkQX5Fo6ZnIKrnxR2I7y
BsA34ed67uPuIuG8aeNKo85hZPavWPYfyUAllhTv9d7lLiK95wbnZM0jTSKP
Q8om3UkXrFjURpB4Nio4RdAGLQx8zOWRfoSZXz1msWxTZ4iHqn90C9bnanIr
95RJlnbxuoyTH0axFe8mOP+0N0sUhWAjc++oIwiRAHzTM4uEaMwxYRQyAMyC
ii0GjsLcUMwMkm7ilxXM5RXSEXqEbGt812QIA4y86vJx6Nlqhj+Ustax1KC+
AQm2U/Xs3OZm5+VsaQS6oN/Xhh6ftB1QJ9Vl5dhd25OwKI6t8Cspx8k264VU
HROC36Fo6zQMpa4ZokPm8pc+q9Z4BFMCzeaV8xAf8GwggqFp1p275VPfLlCu
yDUgK3jfzdGXg+lI3QyZ6EsqTNN24kL3OX94vplKFF2C/v4QzkI5DSzBb7H6
pwTJyyyXOAtvc18bSsW/bXK664xPKx01gQGeWsgmumM/BqONYVUl9iahq1JP
JwYyQjA6RKME+GBQnR85cR0UlRyLXrkpIpjspPk33yMzZxYoGyaod2CmV9dj
CLunbVVbXv3UdUQ5APWj0PZm99BhDl+P4TsjGMc5V2SUHLrvarLnrdJ1kJRv
WvctuZAr2TVG94QU+oYNPysAjIAeaHoZp499j9JMf3VhyU+V4cwvCKNCyq+K
sDEdDrpEbxRY49dY6bl5KPsmkkWDaenCAjBzVC82flU5Ab39kjHiE8ZgzF14
BBcoWgg/XQpXMrng3ScgoI1oWYf12sQRcrosoqI7DfUBXMm0D3FbOPCSPmHB
KEgeOzOYPep7kCn6n7I0FIpLCb4PLdvOChcl9TxIMqpIgIYYkzWE11DtgbRE
PnE8KRSjSHrSSAfi9Zw7H3i0DUJG+dh0vNw0MzVPA4O1L39gn2yasCDwRnmu
3fY0PBQoIKRrHgkCTLLmB4LiVuAiLodvUtjTtBzbuzci/c/uhXgl5o/OQ/JU
d641uAHpslrcTx+HPU0Ow0wWrqs6OlMzfEtyVwpBvhyDLVwKs3GWHcAx0oGJ
FByw3wDxq54oF25Jjz9IEK8emihoHAZws257zpjYuVTZFoWm9bX3CQMmYdbq
kezrZh4vk2iUA61QqWqHXDp9JBqD3sVAc+vVkQCNZxxylmLDTz9vFSc8Y3mv
TsaSnnMnpLEpvpvU+I9w3G0NL8C1elhoSp1qCi+J0F0oRhddDcKtjY05ATpV
X9sd7tmDyZJNRa60ics/o2cBUtmB87BALMKbLY4r+a2vah0FwOXh5NqI61oB
upQuy53HkFnD7giqXYRJ8ML4VwqFD2ugUSG9EpmIuX/VVfcSZ2MhVa0h1FQW
8m/JKsta8Z37Xg+2tpTHOuCakLqvmixMLbJ+tfPtJKgXuc5MLBQD0zNE4E/f
VifbWKoxh98a0+scpi3Ewl7ZXcjEXucMJif6bYbgC0Rtj12Nwc/suP3xhS0C
jw427XoCnLzJg77T9rhaZgfy4TkgcZEXkoOIy35XaIGToLLcYEhWD4KkfQq5
2HY8/xYASDOxKIpCn5OWH7NCT7SWjk5iiw2t0Q4avtUPGcvxV5LV+C72Gu7F
YnQDZ8ZpF3bhX9gX03iSkmkhxXj59k7tQW87uzKceds4nAlTaO6i6qejc6wr
1c/E4t3ypn5wyJdE7D64eUKnKpc6D9BSeG8j+T/NTLeHCPi5lbcxxkiz2zzM
MpUsDTKdW2Vk70dCYXIyL1vl6qOekaDL3j3zG+pdZNlqWXlbwfKfy/WS9Bwu
RBBicK6uiEJ5J3bMOxDgwTUAuDnigbQqkVp5ctogr++OUZHVKaoIt9QdKd1r
4tTGXuMyr8zHVP2rDugLCqdsvZDYfk7KYAYc1ql8ytEjG3dHDAWOja7ld+sM
tG4UWdTtwNSGp63LOqcJcx2iL4kNxxOxFWhDCvFyfhzo/ct3dZaNDPmR63E1
0L84lSNspsBPQKRKXWlJX9qgmTwLKFR8KA6JVw8H2GOzr9eBH4fTxsnPHa1Q
DUD2YLTdcL2EpOVUXinnLwWV5vlfOwKNoxXi1rcTBzHk+S3piH6DZVzcDxr4
qAjtPSZWsOtVo+BNt3GFnWfhwWAc5qhChtMs8RMc1iYoPI+Ky3vxgjSqmdwE
htmCJD+OdDMpx3vqRaLGyZmFUTs8ZgPbWz9CqQQ1zoa4qCFy1b7/NMw17UrQ
sxDzz2jX7tecwWFSnfcIzrf6a9xDJ+jm6OOjJ46fY6EM4jvEJZDx5fGobXje
4GayOgt8cbcLovPYeeJJOGY9FbyKYQ1Za1Zl/nemSXRKa7sXOZYikODn4BSs
zmkKmEzAXhlVEqsAOm5by6b6VWyRxirWYgdtZn8V4uCW82IjBf6bh5hfn8KY
9llRbu4+jRH9vh4wnA+TLGnTad1eA7wQQy9vFMKO72PsWZBXZ//kwAQLyPZj
2Ivcet8JKhbbXVF1+h5DeVPhlYuZaIMbTdIEfHZspi2TY8P/HLOV1mxKsaT3
F15f3XhGDl/EdCdVeAddaPpJUXyog6pBYJFINjCFef73uM9CwA/60kg5hJKN
cUGaG4rFBaamhvBkw/d6avSeJqoaUm9sLfYq4hhzkulDwCNTMBQii9JRBw3y
+3ll3a1e6/Ogh5O39KyIoDpATIiBt//IkS8i043lB05E6KJDHtbOv/zQmT5x
kDyNAWu1/hltM/PWJXvQCZkp37OoBWMztgGJapF45ORQAIV5PTYglcxheUp3
i3/fKGwdGlGvAe7lCh7dgdTFD2iufl6wUwl1c0A10TzsyFQc4fiGCIID3EvC
X6rPZhRNotO2jGUAc/YgzXZ0ST7uPvpSrqap+7sV4vi7QEF1JC5nVFqZN/iS
g6u2ZDGFiqerJMOuum0yqiGGZTh7biPsKfbROWhRFcoNVMgPdxOZXhYLvCoL
6R91r2ZepCt33YNCyAcNwIx2pP5N2fbR7UJBoYBDe60vwpO/E7JlXeOve2yi
V8/T9Ll4U3NShhK1ahI57X2td3AfRLBlF60l25AlrZhqzqBBnNBgFGbnc5xs
a/mGXKBE/Rcf3fjfUOn4urqLxiALcmtTPxWgVWK1LjAg3+Nmi1mj/gHslh9k
GRzM+9VxA9Pakio78JGJObc20w/9VIel/tdWVFBnHjEtnf7zrARlreXwQr1K
0SKsb5ltlN2rPuSCw1rPLLoDvXOZq7HRR0xxqJeCxYlbr7MAx2kKvz46QOdb
mFm1Tvr5nhONkKHXAw4np3gO0uS9grP5TJWneXgpgVtbxNZn+T47k7olvUnE
QO8mR42AuVrOK1qg0jSm22rq/DfzEoClDJ+Z+OXzhAjQSB5nvBosXGB2Yml1
jkuvzL9NYg+2tLPu4XtLhISM4azfyLkEjrIMdcdWN+SQD3GPgvYfVuJHsBhm
m4uIQfKSg6tVJDTs/JBTPlK4NgtYt9KmRRWjqHTzbS2FUuhyV+AaKhqWlMNd
BqPFf9XRACdIdyppqABLoRSNkN1sIYwcCQzxiZyIpCO3cufP842FPmKTqrRe
tt4bgIBI4fo1Mokjval3waVDFlOAzCW49+I0OriY1pd1AXEf1H6XlWpT6V1C
jXc0mHENNXhIcGbRYkfP+6Rd3nDNEMqyP4Y8gHoVrY0UDjENxeZ4UdxZIUvO
qyyq68Lc0zgYTrzx+SxjITXUGNHiQZAdmmT10a8r+HdIxeKxLVT42HBjz89u
jRFdVjnfv25dbPk7Na/2q1WNrr4aK7nijfEeAnBkV9pZYnxvkrSQCF2ER8Fo
41oiSq+kJYUGADsY6ETHm7K2oy/7n7PJTkvOzAWuCpWonf7KLD6N6V5uWqj3
GIL6eUjV0XkX/Jw69IyOboXWScVSYpw499eO8ixSPe9uW9mJT/oIEY1YVJQo
L2lgqQrs6zITorOBKa2qy7ojhrko4t/jeu5ZkNP1V+ZB2H+MjnhFIElRYi+X
WepPz7WGe2jDtYWElsquhgFyepnScq/Lr2Ws1wkv5YzZo45+gHXMqHr25g6O
+5NgGI3L1NMJtjP05mQAUsL26vlbXRtGcl4UG+/E6rNDQGAWod2GobMDUqf0
kLD8SIn13bVWQeXxate3DDDSI5DFeaW5cprTDDqofbgec0rbi123ffUJOYR/
4BQLEO6JYV89A9NoAZFNlHI3EP3A2z8bFw0NS9hHA4mI+Z7+cDco2ZaASwRd
LkCFVDz85EGWmBxlfRIrq2O8F2YOJdSm4NikKiRoJ2VMKaexqQCC1hOIah2w
i0SRH9ZKxP+/ymm2uIIBX7ZMjDD7FBLgiW2E/z7ynATIMeSiSqyyFgrbgGEF
+m2kGUilOLy1FhP35Jw8u/y22atLvA2de0fltK3Xq0q59Gvllk/crBY/7v3H
qDH2xFPHLDQQBZlST8K/UVuXBeDqe5+rj1UjP8YK/MtNCndaiNtafXiCrbK4
lVTK0Fh7zmdhcg7LCJgmY0SwxiGoH5wl6GKVfUQzK7tD4bQFLvA2DmSuxRfq
jCyHHed2be9gNknos12zCpAXSo+HfXIJXBq/RXN90eABcCsyAOWDV15T10u0
IMsQ00VcVyAaQgBPMXoSadhtcEAvo3WgmVHu/G0fX8T+BLUUNBEzyDe0pbRo
EF2kDjWu+H0GJCfh26ytmC61j0/0aAF4OwdP9ZqUyqrV6IVXJvXJNcfitPhc
AgcLrE+74Xvv5APsTocteyXuNNIb6RPa/FEVhsaUNW0ragvhNqA4WPCV1LmG
bPJoGO4cxfEvwf7/Y9zN+D362aL7PU64ZwNBp1e53trbqgOVaBVpv1Qy4RL5
XKZz3/rhLJKwXmASihM7A0WbqIkp2Ss4rXvSPXsT7tTpPY1uTKG0grwH3ZLc
sV+xPClTjn9i2T3GUKlTY7JW7+F6GLo6uxFnf3EB1e+EO313bODABJdK4Uf7
5eR9hzCXIqasuX0KNRPIsR5699vfFDzfL41O0kkSlSygkhTu2hxCpqQ6neSq
9jYvgClHmmsJ8OvB3y3cCQMsoCZDvj6DFHAw2d6Too07wMe4S2S32i/tTGOc
sPtsTmvDYNMyF6a0UddAWxLYw4nsLOP2xRFjaHb7F4lFpnhvNCCtzOS4PQb4
dl5gBlBAA3uR74EBKLmRVBgsNjfFFxMvFcNquC3eUsgX4fsE/0WpOig3NLp7
rugyuIVTJyGSFNZAJceYQHiUh0aZTse7dELw86UI1Fqcqi1PeZwTrQ/R4wVG
EPEP81oV7nF2trFcKsju71UY+5H7f32P9yPH6o6Mk49/kcGasXnWAtUSpg2p
u2s+4/fZUXSfS6rnxIj16MB/xCOGwEDwN+Y77aLUkA5AjjvngyCjLJSRVh4e
tFWznc0Zvrk++VlsGbYtSWsVq7Oy5tcWATEWXn0UE1nBKdnoZw2IV2xwDKAC
ALff8c59DlYa5nfBsa+OLDHNZfUgzit/RKPiE/r8qQ317OpKn7iidc/pyUZz
PTd7ulqS9CBs3jIgBeZlpZgHFFsVsmuFwCFxZr9YzWSiXZ90f0cl7lbselNe
+FPQUHd7rCoD66NH7ByyeuvH0hn5ure8SJxnzJ5lmxih8d3IOVukK8202RwG
OIP2aaTpZlYsx2I2u5YYJo4gemJ2kNkbAC941cA9L8RQwK7rnh7XWLLY6WrN
uWD1deW0ixjOktJqowXrSFNbeAUi3wlFEkv1NcC/l57IhgkvTNIPTBxRX8vH
cNUcXICSFMn2yrBJzfGTHdJXvCFJomFlFJt5iDmL1YBRejU7hGZqJC9EnG/A
cwZikUc0RrF9zp5HTvaNaS3eGVf5FZMIZ7t0uI7j1bzlNUsPASuIerGFE0oA
vq2/avbyOL++Tuy4QQdRTpv3IkO1ImqtxZ3lz+OoiwNRJCPIXLYNVdQtexNi
uWtFZAJ/alVjlvQYkMPqkt6v7BjNF4b2+xr3X7mQxgaWBKctandJMMcFYdMY
RDptggTB0LQII8qjSIs6JE7fI949ZGsPKpxFoMKF/N4+hdhhpqeEGsst2bV0
cL7PByPgfLbZITYOLbEu/pLMVayAV+u+wmdU29gA35K2Q1bre6E3EtsMYqox
VmhPi5CeYWFd9ikn7B+Jes5TAK8w+EC1Xz84j6Qq+oqhSXvwHP9KxhuQcs7r
66T51qUuPYcjLIufudqoq6Eg+olnle2UkfmKSl8w2xa+vX019dBEPu83+aEw
Sbl/IAr4IPCiJszwUJWSAXCPgTVERxeo1hgaTVEe9EqfcwWg5/4O5F+RI7gF
zXvkmGqBJ07GL2zkXO9YWhlpo0dGtSJqnV1nlB/RRvuqtBoanxU3W84VEfC8
Sqz+PG/sj5SteFHWwUK5wycL7AQigAwRqbtBvOHploYajfP38YLUJkAvbA8x
3550Wx2n8vzgmtgOxlVY1+mdutAi3YGdZX/F5bCQTkTjNH2j0QhsQGugioN6
IvzIdr70TxcdeGx/q64VOwkAiQW3zqm4osEvY4Vwl3X2fz52ogltDiEpD/Vd
Sb29AvcDD9/w48KFoNPF0O/yCRBbOizxWjwgJTVTAwNbkwCMhizwJaTKB5E9
WLOYmpAFSR+CrFjZwobN0uYzb4EYSsaSJQ3HrklBgDnFHZizmfNIpqWQlnEW
D8EE7xSys/YUfHlCB60DwJMDClDbbdfbKgBFvARcXOJ+bHiTekr/VH/eBARE
8oMwJpfa+XbJI7PipTtNYhjHWdv9XF4MzrwMNM9MEZfeuGFVmZ3DC3bPpnLN
IZG18h17amGpBuCcqMed1RksD0LYxfq/Pr3/smrR45FpRVKH52P4o2brBtM+
oBSQjCZ7DsIlnAdn7xYFvX6eQmGIkNRT2Wc/iWRmPw/ELz8nsdtNJwR53lov
HeDquhLDl/H1e0MQgkXxEQQLtXLoH1XeSRQJyKcNhKK8lfEHvDe4Cf9OPPbZ
62A9g4xKay6tmWmkTNA1YkdG5rN7y5nilU4kBsliIa2qI9ewKsAXlrO+VjI1
62brmv2vpFM3b8pDEfmeM+CuwEogCb8qUVbdTEyqT9SgPzHei/anIed7d3wb
bIy9UfX/JJ4p1N23JqRNKVkPwoH4xdqMVL+w83gLuMfgnQ/tHkCZxgD1rWeK
rU22Z4T7jiM+jWBuclMekziOEtblDBKDPo0ZSyHxm2jiJYseV8s50FSghVYd
GhDw2wNjEfvg7kdeSZ5j27RGtunpy1lIjptfMot/mglQATS58tfvMAkYb6wa
zfoNUo1I5RWR61+jt8iuNUWQYETn5TAbpxNE5q58Pkg0mFk79+8IlmjmNQ6O
3nc64cywAeOyriUtZ42Ried3ouR9QIs1a0WnW/GoCf0IB11bn6tN9wYIthed
4Fj4R0nF9C4YSfwDBStGam3tYYU2xStw7Yy8gFvpoQc3W8i9BvKFAyTtn+ky
wEjX6WTIakB8HOiQ6VYbU8c52s0IkqtZn/xpKZUwTunk5qBEcB2sEashKLin
b1iTgjowApVFMaX+vqec42B3N8nDyAleNOtjzkVhFjr14bHDjPPA+t7Y0yni
im5mTT1xwqfCxOeb53wHeZjZkVHAqsBwrK17VXr3khbASzpKbo44zrwIl1S5
k7WY9SUKpvi0MgPeEcZ3OM6szgf1caKl+mCM9G3HcAYOLDU8ALLz/3pak19N
wzjQoUB8Aojg9wB/vRVNHtW3TKLiaATnMDMCv7wwGxCsGKJUpO4I3pKO6jlC
XDLSFDrvUrtQJ1EmD4SxmeUdLR3VfifWhW3lucosCzikf3CA7iOn0IARTsCM
qU0bYPP0N9uwMrFRzowaeZ9dSRP+BuYaIbBxISGvXvBcOurpVZUdTHBQJlN+
qmnlV9G42nbaoVJFlbT4UXM0t7XYJM+eUJaDUeKfEF7TTPVQVGEBZBGDrAAd
Ev573TbzhvjyRy0WTX+ZKKMMOt/nFRFfqg3YirjTL0fvzbz2Xf+uojpJ7Kl2
XA888z5yu3jJ0sNK5k5JKfKsBkL8wbuFsc2rM3O+XM2H0nmphzUDeGt+qcfz
cUaK0O21nsIRerkXr4cCUPcvijK9E6HGe/6b0/3GvxvYSkcZ+bW7bT09uVI+
L3/UZr4UNj5/ki0zvSNO/3IrexWud1EkxI3BpiSy1Y1heOksPeuDm18Y5GtU
2JKO8nrN9c+fxqlVq17XmoFE5VgBdS9lFZEVovYhGb4XxXA7lK7+NkbbGOhs
NQr+HLbYtaw1E+F3Zbhx/NFIaPC3N3uoFYSnYezaHVc0gNRkFOITP49mLFHg
nECRHD7CoW3myADgmMwurlp05XhRCFHcGxyebVgBRmooEaUU8R4Ho1++1Blh
szNW5268GOMb7p/9R3XFotUBoqwy3pEY/TChetjOeGtfTir2EkAl5RaxPE+N
kvolHAOQx4FZHVRz9a7D4i7bMJVh3Kvv21Hyu/FVFp/xZDY+P2bbdmlXAk3T
NMtHbV1dFA4vFQuKopygsUW7+UhXSknxXS8lvo75SZVms+V0T4O0l8H+51u7
fDljkadM3rCfpPnSZ8CHeddgRGB1oeyDk7n3pN0Swl/2CV353FyaqaWQz7E1
bW6pFSOmvlukM1WMjdajn6lYCZ3wkzLopbYJMxSmPnhm0nWz9FG65y072pDc
TGUUjNMfpfSt/pD7n1LyThiVsHm9qhyxianQhZvrxX2IjnjwkAu7/x0DPG12
3FCk2jTfh+SJvgPitTMz7NwAmprUC11AlU3mCmHZ0zZw9/r28UxaYSvYS/JX
/d88VNAlWQeUV5Ph2LDOEsLTucdjuKCd3oZAPq1J0/9uQc8iAexjw0a9cuoo
myInt6ObY+m1BWjr1VQEP9jXAzsu6MI3M/UGstvVQXtkdVj8ypGAGkcbr4a3
aecJ2ksiKmmQGrMIZB90i5LFSdcjRI9qz9K29nk/Y8mzkFO1X7wusQ4GrfbF
tiYG4tZh+h2RgGjXNPCwumqFgCJUmpNBq02/R1UGFjEMULpQ1mNv0kPmw22Y
0jXIusTojQcpAfZGTrvayWkegsSU81JuiufCjxJNFbIqXfBk/ZoAPX/CVAGu
M4bJrfBXbfzUqU7RhpNLWI9riyCaVcB9g1hSXLWr2kBFFR/4b2tWskgzxWfM
frlpG/2QEfQ4Zb/q3T+KyoetJ2dQatHeja1jN5uELc3zDLKMxgiRfVfl6M+h
2HzX2hUE8qT5oVBTiQYrPtDdCPi3LV3rMNhDa6aVeVQ5aog80czvLW7W3MWp
Z6+1pidbS9muB/qMimbRP74+rml9PMguSaeY7Udp+9n12LLZ23XWNwuJVUOE
HIJdcJi62l2cV617orNvD3f7WHeQrPElqKYDwowwIcaUCErDsV7AjRyWpIEv
4D414MCwCfR0RbMi05lKDAZyFIRSKIpey2YboGly0olUqDj/q3aN6Ul5ZpAd
Hdzg5BwUl7ZZ+TVrtBvdK7GAoiAW3JhgByqJ6UAjzJY0GibVsPDrMoij58YO
EVuV8bahHfrjIRP3gw7B8+/ShRwN6t5uVrpfs/ySmT2c5aTFP8tzcgZUAmZx
zH8vXm1WMF/JUvGIM+mmvIc9ALTrNsqPFOBhDs98dQVCiv2/a7wYyhvLVIP0
XMBJ6k1H6t+k6h4EWWqGEkiqkEZDF/rMNHIJe+uoWHqi9XCWLRuxNsHQdCXr
P5Th3rhTF/Ibu5wCadQ1OMtJTteLQ6s9oZ6gifjKJtoJkW6ALON8MKDqMrxh
r1tHwpJ+96bwMVIVqaPoHV1BbucEVP5p4WjW97/U+18f2Bv24IueiK1yKSQB
Hgg95wPSWBq5nOC5vWBvHnkhMZnSjkWMO2wOZUof3E/2uvxSTpnZUkOn5oIp
07rByT278e+LZI+G6YrOJqvyrzLNFyHEEoKLSFcIw96W8a9eYN4ro1A1jind
M/bfTTsXfJqUWHzb3RQjOmUWUALRAzdluuLPyxkgA0GpWbmgJ1SlKT6p0DV4
mlLVqEPCNI4vrHN0HcR0n1ycFXuTJ/I5I/pDyQ82OedCJvuBhsI/9pDNve13
fQvgxr/ujwi96UE8tRFqMH7i3maIGGRu91o3OCHenKBoBWGUN6s36sB4tkhr
QjV8xpkKFqcSzuE4S/FYgvIZDJ6VVWmy/aVved3msjmeQh+/ROZgie4LJPE5
BhbuovrnLH65EzwAufrTdDaBcWQzE02Jo3B4ho2DHehgxwiTYFS+0Q8PuoH6
9IUONlFyvpEICJcbyKB7EsErgSOHbc+aIvtdLkSYLb2Fu3DwqdzQr4Rv1Fja
IE+xC92R1lQHmuvN+0m/reAUUgRey6szQi5PMfbikrB8kOFWQ5y8TD0nA6YN
hDO25sxGBLhwjVrutp0KG9y98ESB5XEU5Gz5tN0HPwGpLrJnin3mDQe128dv
D47VYdwZzcRQgsbXb1uns2SCu8GvTVM4pRnuwK2gfwY+lzEja6XCISiaczep
LcKq2MT8uQTOObLJ54KoXyg+syP69tlad4A/zsWi4ZeAMOnqS7DC7RGt0eDz
n+jKvNC1FzW1oUyDV3lqiQuqta3o1M5QyNDSxKlbwARLVT5Po3k76l965oNQ
AOGaIxBxrpVCwqReqo24Oir/MzEsIz2oG222Zwm5xMaowreERrPvYUBUDXZ1
gNOAekVjQD+S5Kad6dRJICUoA9O2T/AVVQTX5UeLamOsSYACezMhWMJSKHGy
Mted8UZTCzDWTpcsMpunp2tYkPjmWORwq0xMptAv0y1aEU4CSnXPdY5Rb2IR
PUCnIbXLPBdsUEaZr/83cb8+kbYDY2pHsGUtEnj6dmbbXcx1w1NUvZPfCBkr
xaqhILOtuXBmpEFpWKkmODWhqCMHuPBwm6Rl6rAiY8+62ueO16Sn1tPgSqaO
PZvuuW+x1X/iL5/vuzhy+7vwcH0FWSzlMkMk9tfJRQs1RaEIkTme4yYJ2nbD
eJMH/fKg2sNiULQKmm84yRCp8Ha1/MnzOXQDuRolqjT8aCxrLdAV9vKjdkZD
013RrEMdUJHSFoxWLVoDaDm4HRJI7wp571Q3lBn5GK4KszE0wsXjp2IA/Zp5
xaX6edxlAXCO5ywKyTuocF4lHrz7svvWAPrRupyyNOuRn6hsYfR3JVsRnz52
VrkDZfkup4qjt5XEA4R13VqQGRHmKeG0o2y1YJuWcBijRitzG6YmyVjnqsla
wvvRVUWEpgbxPGxH4S7NG/EQNt4noW9+8LoZnDNrma6oaWX8YwlVlRbuXZNA
s2V/R1f0hAJHCuy6NvgsHmPnHNUI9rMkgpwCbRHf0q5xGBgNtkW+Y6QKsrmq
SjyvqtK/vRhW7J1p7M6jUDOMkFmasaK1sDa0

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "q5w9/+5Kue/STKa5XRRpVGZJHL0ZJeEz5bcA85thYUmp1PIQq+G78CEzW7wlYTXVo+w4BCHd3aSh/18cFjiZbvt4xJJC7ehpF3+ycjY5Nbab8XuVBxV0GtSWyUB3OY5g1z7jhNv9saTklZfq4NIuPRMvUINOi1jN2p9Hk4oe71H1u1YzS2f8oWdLZgHwWW1RhshdKbt99NlJ2sTPdlYrRV4HfVHdWgZ2gEOhvkVbm0twMoLcB6cTljrVYfnxLPWQ+C6OVzbvSTvPPXeFd0Oymu1mripOpXSNKfXOqx/wfJPL3ZI0BTWYEeCUUv+xOZLbWk/bfUHug1SNaMGpxom/HR/Xf1tLAdjguvLFh4QPwK+vBUysd+OFXvamt3QyofCIVd4kJSHn3rv+vJ2j9E4MEldatQ9GFV2pP5ttob1onE6BjHvHOiWB3D+YIlQe0TMqyYjmrODCnRSs9mKfm49RDqtl/m4SzYhyXWq9Rt4PJS3cdzaqtpIqAX3rh4OtHgb21oDSr6NzCmbLhdjivBW/P4AwN8KIM9fv/qRePGwJAx3ijsGPppDoohNgj8e3NOUEd3aD43yg1vOoDkjN/USnTGX2e2G9+RuZbBBt4pPGVwHr5CllQnnXME78foiEKO+xg39D0vNToGvETqeMn5c3B4RXuoNgkPeflAJ5+6vTkaeFckTR5C+0carek+rCjh9dK7k30y7xLWtJtg4HN0E86/a5Gqwu9fSFm4UtHQXclpwSnkjUFAPSEdjCsJZ62P92xSO2CxQrYryl7E/AZIvI39CmDfun5VE5dD4v+IWNSUjI70K2EFv0n1FH7NI1Tl5EzMyqL9v/1yA36mSzxPnhtHMIwqRcTy0YLYdc1nVePZ82cnD6h/XUFYe1+JKImVtBeI0GHwOdcfFc6DHmE+wpInkfofunqU3dIxY5C8LQAGbLTOaNjazWXG0zC5kdnkfI+GQddKqNL96rtIu7R0Sudx3XfoaOK7hDQldmL3PE/EDfoThtBcbtcUCYRvsiD8Cd"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
btyaCE7fh6b/3R93xeO9sPm0D++z0F6iygDxCVryt4mkxEgR8UAW+W1HDwsi
oe/rQAlZeuqinwi6R9tXMS8keCzHPGuApq9puyprM8kHXC0vmD0ndiuWGJIK
y7VrZ5yLs+19ryaT2aNkEB/5pEfhrnfisXeTwODJQNZ00sHBV6bLhiIbIO8H
WKMJ6vXSCcTJxSxYkNFlLR+fIsJ+4ZzE0U/Bk51ow7vqVIw2CyZ/Xh6MEP2V
4VY/pvOsyKU0m7hVxAqXxPDdoNZRIiBjVsb8F6bszt3LNmPmBlxSTAZFI9J1
b2gmdR8wOwCUexgoQUDN9tOiE0qfwc4IgOZ7vtCMFA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZziVNkShgBt9tJMBQXoU4ZIDcNG7RSr46xACIVTCm1GTjXLYyYp+6Koy0yw5
ruoNfICVS15Vegx9+Tq2PE3GXZhql2g0lcOfjHbUdvSwnhwq8aCnYtR/nY6n
O0VWvzSjsXMRjSdnR9HaxjuEUOKV/Ez7RfrELEBrY4kWdxcWbTNNPpAKf4au
Z/8rCb4gk0/jLrz8t7Y7lzEPEVXOX44RMTR39q/48rjXtczILOkkQvX6OHFa
DgKNfiF3HSSMedoHzIr6qhdUNCcpz1uUgy9ujGHZxhGPu+J1BucJN1IIabWj
w5qTNnvhyKHVNY1qTTj1eibY1flcgKTEpg4Q2isTEA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cNdiaMObs+6HbP3hHQwobT2h+PB4rUh/pNTGsgNJLhdModGOeEkaZs5LHjXj
9glBvljMpqIzbOc4B6Tmqi+5MGmXSH4Su+AlJFALYy8q7OVt/ouZm1PAX/OR
+SG0KiRQpLvJhnl73hV/Qwz/cTHW3U+CxDCn/v33IDyrWrRM1N50UGz9vuRQ
nvkRW7OFY/Dm2oY48lw4zcAWLHR5q+SuAdx9YVQc/calLgk04JoH4recXCG9
aqe+Cn645bbORBbJ+yKTKPatfM6XuNOrt92rMWWhImyev3+vea7ktmk05KWG
P9mbV96pbij0U4RL7pGuTKmmWpD2u+hyAiNEkrDRnw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BLHtlT+jTWKnl7us9hBix3Q3C1P8TV2fGSmIjQGfhDWCtA3n3rhQmLe26P8K
QNPR7z4KXzsFl7TmSC4RUfSsBSnvNert0+K612HKA3EMkdepeswr00RUgMy7
/V4yayX658dr1/YXTBAhRu8ye2/D0z7gP8UYbXK1j2SsL3SKKOXN9+D0N1y1
Zn7Zf0fHUIyoI6XBJxHlATxwa4qpFe8GGxQ/eLbvb9FU640A5/SZijSCA30y
OVwqJQvVu/pMhdTV4U4xxOhWgHF7l8GRPeTrfu2tbML3zpE4AQDH4HAuxL/I
5RaTb6UXeMckZ/4n85JSMJrCTAbjTJd+eEdfN6aMCw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HPho1HTQe87wJuBqYt0OC9IdEal794HBzkDSkZHriB4+KLydn00CazYIMXs3
+9ZVigUBPOow64uyD3noKiOK+BMlIirF4RkoxvNAmDcz1Z4PV+SNqJWN+kTF
NkgmkS5ZKk9fSe0zcMn634RhSiy7eNRMca26Puzs9wAJfgPRfvo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JvfLWijvV8DXJZIXLIDWjsI3NJwAlchk/gzGI9AmscxHWBDeSNFoDjRjv+TF
bDhui5nPRKNtv+nl33JY+8pFxWyYCGwH4KPfqMRXRbuVYiUKMhQKzWn2rhRD
XJD/Nd9aeBEb2dcp/KmeRTumrDcZbwKGgl90xRMpkf0zJwslsvZpMz5e82CX
CddCLDcVQqyUihatkSDMr6c2c1dXft52ud6cggCjFWmTGRcXLzj9emz+8VUF
IqqN+GLTLMZo+L09b8Hh4tJC8Ft8MdJFX0BwOkdq0D2o9A0Gdmg90i0g/wlo
x8opIMbfraunODn0TOpgebS/cHlOCNsgsF1Zj+7py31mBX4JMO0PaNL2rKnk
CS4z2jEKG58c/g8z0A6/YWSUFgmgR5sjQ0mEZTYX9JddwPqcy7OrnO7cm8Qu
1yR2IAv0k4kpwEjfkHiHyibrAPROdI+YCNDJ5Y0p42Ql2EGZtNvidR6eNfBf
vdjgYhwqCohsLqf9vd2Tr07gVnR3ODu5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Gw+g8YD6UeMmZcMVUj9FwVQsJT0M5bIhIcfR1XRIASXnTzCeyaUVSD6shq9j
r5X9qqkJOqqfb+ebra+V7E4kLB8Iij9po98EEMWQ49ekqLxJuA9y97Ehxlh0
mtyS4RUwQirrkNgBNGVuigiYd4VK/xg8GWQr5/ObyBSIpY1jFUk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Yjh43Psb1BkP6xikAehj0hAm0dehIqMgd/CWl7ZwSRKYmY/6JjTj9oK8feq0
bXKJZ60qsrCSEDvgZqi+ruknmOB7LhM3j7a460CwGou03DUnPiYO/1P78uJN
KtX4KIBwAjpCvLpMcbCHJQZgDvmUgfyYlzXpB1AoJrhECi9yubs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26912)
`pragma protect data_block
/jlBHsO7sA8HBERlg5H1F688RsoFv3BQ6Ok8IfbSLW3ntP0jV7qK5JpK9kmk
2YgLPVgf0QQ5Fmtya78DwuuqXWO/1evwvgOgsdLnfgwRSqQyXjYI8eLs6r7f
XJCUwvlQUY2aPmfvfl6F8gyGDq/HhV+TdyEKp5qshdlMKxXdc2f0JHaPLy5r
HYHuAlGbtobNYUMyogV+hyvwSJOOk+sxxbnioK+MR3JRhC9d88V1OefkYf1t
Bw8kJVa1pj2sfg5PAvC6qyDfJvC5PkpTQdMdAI2ug7EmW3yW6t9OLVbU4fhm
JLerKIe4deSosxPpRtNqWsJvtrWU06XpDJ/MqF0TeJ0eiWSCnuqY+lqBNLWn
/FtIvWGikcl42z67ONY7hmnT2H7qKBMKyA1HkXPlxz6545/Iq4lXllEeWKhE
t8klR38aXiJ3COBBmXuah6oUPnfHbOAJtRvfyXlWl+gnuwMAahYYgjvEhzgd
rW6OzBdBkNMpOw0I0NXO7dQAUyYIsbdARR04cZpf88alRIykZOiqcIDAJCjA
2QJeTfVPJi6jvTcxLdUiaY4K8fK9DX36Th2VQyp/w4D4hiqgtZVZcyY6POfl
YdiDuPpgvWbFzvjBhCpuHMomgCkB6dPkjgt3hkw5ZGLA6RG3gFt+QGKKt3aP
ZrMBviUflXl1AEaO0XhAwYi7qRDr721cPBQ6oCri6TXFwSTgK7lLk5lJUtXC
C1XC8MxGtPkuIMWIimqoiA5UK4FzUy/ZJrYzr35SRBzJpRMykavLb2XJqwH8
LiPcD7vmXH5qnhHeNKD/jt/hHRwdYykE/Mpg/X8ktpkO6fSSPPYMehdKq+ih
oalzCwY6+bKOY8Lyw0OCiep5vSRJwqIrSxPIa50hJjL6bu6O++Np8iKQHP45
dz6SXzB+6ZNr5hIus3zIWF3VlFB5q+9qJP0sgr9fo/aoUj0yVLidn0kNuRjL
9l4it5k1cyfpyM7hZWsfi/0aGRd6uPJB0baMmpFxfVeFlTfbombebZ6t5TKK
83d7JzLxZcdbRbIhxgF82ZL9D/mTTR6Rjrt89gUd0BA+azxqt+w2JMejYAgx
1vk0b0FtkReLynxPdTnz/AgbzwlVGa1GQVZBytgGe5Z7uEY0jU0CIrtvektG
rg+JvvuBfLWMala/3oOyVHy40VSBgOjO2ioqc/B5dTKXmPPtBj+sPqtbWkQz
b+pjmYGBcJ6mxviRwl6S9rzmgbZiRnuM3uR6mqNz/Ly7g/1pGvwBQ9ug6NwW
4xpQf3vVqBsY0+sJgvSZ7Mf19iyIj3OYZMPfA6Mj6ga7wZUAB68T3yKV7+3V
BTniAFcopHuK/7sdkCK5iU6nrm8gi+E4y826BQ4jFoVvorqIq2CGsZznh+Xc
+Yk0DQDd1Ndn1YSdErJGFyEpCjj0OZWj2lkFU3f3eAfFcAbjI+sdYwU/AQFh
wl3Bbfll8g1h3R/LVSCUgz70mEVLbxOSwn9OhN0OueisVqYOKMXoh8oYAvQ7
uNNfRS7iVKAPNmKeQXXuKNqocqxN2Z6I/7MWtqgqswd3FuHNp3nzstXrjP4V
68LeQSw+eJsKrxs1EM6m7is/GuhPzu/CuCITQV8WJ45TB1mXFigYMv19g11g
9ODD5EgosTociwOTtBChdo008Q7KGvyhVkp9ddzFFVz/FxCEhMhtRVtL3v+o
hArGusLOdDIwaVE/E1+Jwx92S8/yEk07Qz1oFkSmK0xPRvoJmrBJMH712ZE7
D5RluP5n3X3kAAFw3DwWY2JS0+38UxYKIzZN+nYUBQCZxhxRH+QgM+5BKT//
JGenwgg1mxVYDQEsDsqHE8neSmOSSotum20IEUk8HD/pQaZE2RJxib2EvLob
BVb+bdrP8dgP0snMA9UJhlMO79OqtsIv4Xrv0rCI+Yah7o9U2+rXao8uYiY3
zh/7Wa8xd7NsoB6RA+uiQLrUkjTASye6O4R6FySnW/n5FaVuE3ugYs89f7WE
0dEAcJItmsd//XDpVDzDN/lpNsE4zAzKPnfUjQID4fvC6KB0Gjt2vwIpqtZh
phs6o+exTHITDIqUWSEgn6feo9UQcL330kR3gO4JFxCFqvc3OWgYKC42ZA7Y
bQF8EbgVM5BbWQyStNy99XrtqWVb1Z3XiojgOOoOSuc7wj3RPloXzPwZl9aP
jrhciP/a/3li29PKmSnxL3jjG7jJVvi8OZdBhoczQVtg1HsgZKEDdd84/4d4
GABevA9e9h2YsVnlvGOE9fjsXHkrHPlmBUZyfMs0uxmJSyE4NGek6kk8DPIt
c3pjAQsp1mhUd2DL3RZN0mr1HMKESmKz560mDrXird9TMjNAdNRI6DyWn7iG
fI/NrFSVYJzp4WpY5f5nyJ84M2C/DH3WFLuUMvrzHvx9QpF4cspE77Gv373r
qsf8yk79AncogwmfhG4kliqbQKJOB0MXbnskuspr5h8ep4PWGSeY82kxYc3m
5CpUwsniQtMsjYgPAtiJYjbTJmDD6EFez4R36HQs5KmXmug/z4YOrH9j8zQb
K66k88siPRLsHbIMjCu4TBjD2ZAkUMZN4GMxeeOrRbn3UQ6fRTusLaLbpNUY
EHXXIbrazi5aEJHjFby7pdQFtEd4qcX514ib22xK/ZD40COC1ls/cihGJADR
QBDDk25fgX2t0Iijt6VLDC0el10VD0YpwiRXlLAVVtRAmututO8cJAIHAejV
qfY+6MXPNCW416363IHFA0ebUH3l20hU1xEFVkWxpqzgjPG90sNnDV/fErUL
VTIlu2Y5UcTXoYl9mjYPTasQmDifAYWmvjj56gt9AF0LuBkZGrwcnyx7Wi8x
xcCdDO86p/dO7BkdITyUqc6iSHuRVXo41STdOL2+SzqX3o0s+kYGsEvSiODT
UBwS0PZnYZnA0szkv0mhfqUPruotpav1RNIFrcwMqY9NIoWi3IePn+cxZ+Vs
WYIznmwwMV3pky1xU9VNsae4SBrRop1TMyDj9mPDWEWJaEqQQWs1F/RI7PZD
hFu1DdAGAYNlVnOGi4pqTk/60Tbypi+h2yDIX6npdmrfmrbLuFlyVcoz8ion
miIouDhO3B3tQrL7kwqLHveHi1Y+ohXHGYnQknQwVh3LOZ+WHWy0JT7oEVuK
3gXgtz5YpDg98ouTEhg0TsD9f1MxCKGSptWHeKA5Js+hqjtNofewTl1msgGu
Fl7pGCsQycbXqEoY1VcmX3+sYJKA4TxFGS3yBIhekG8FFM/hfnJp2RMv+G7c
q2oMYXUSE2qIPK0GDCh76gW7QD4T5NB8kz4kW9xJbcKAcLFRLM9M+syNowlz
xtiovQX3xJHRTZXbXCgGhS4mBtoKSHJUwMX+t0HvdAQ2LRORp3DcX/w4tJzf
PWbTNcE4zZLkQF5FAN5rkQMPSLUVS0plzhdDB4gFg0kjm0Ao9Lz36BJPv8ph
O7WyUK+8xmntgFTzrnA+F8gKml8emEVzaWXni4Gz/QFbsPC0iaJThaLgNyYm
3/xJziJIQY0sUfS8wYyCUPzZqyRvA1iKrhT9L4bEUI7CsM8cqKUw9cKweXBB
u/a09a237/tfKD6fA6hz3B9oSMZo4BESdYL7Mc4ukJOgg1Dj8AUdFfOXS8Vs
1TaofAYkdriITRswGjG1B3FhIGvwJPMzm05DswO+p0fdIitLxl4A461BsROc
lXOp8qVB+pPid2rs7jM6Rz6YkC1LJaWIkPBCATCHBw61a5rh03AjgNtykE2M
Cy3SPGuLXUFs/cQo44WYrZTOuO7i3/dZGVMSYVr6tBfqD+DCanCPaukKZPbD
PNfYD+TbH0h42HJxg2K3wW1qamCohLkZX+B1Ph6QJ2YPZSjllpDMV/LvpgD4
28sKA/dwzKDx/6fPYpBOGJ3lru+B0rVdX+PO6izLI1QDUDTCea3MAgF81wRW
IYAP+4YlGz1zb9+Coy+wI0s+yjSPG3Ng4pYemQUHw7egIDE8rM34qOk90QXQ
84q++lDhIbyPwiQXamV6hLc2njX+409W771EI//IHaEujGZWSQ5oS8RtDXoS
Q4ZQkrI/39PwDjKDv+P81AWR0kU5jot/xxOFwzRCrbmPe8oM5dzL3vYvGFRJ
nJfkKGHI2jXd01xT+TmzOz0gG9Za6/FCErIKNAOEC9o2is5aCAqImEMESCjx
3tOS0X5tcIS0p0bBa597LZKjIR97PDog0py5WEqXoWUEfVFjnW5DJkh/FLdX
A6Yva7LytIEZNLOS2SvGpb/OwEUiyoQzBTJ6kYk9Wm/+dHYNf+sQK8jVaBAG
vaRYKCtllYpR/NRRrPiwrhrnHC9gdkb6Wk0m+wp5ZZ00Gr26eH8HlYUmBXwq
5EMHiucFJXYH31nA2pLObE8/2vvqf0L9T/VSTlRDFx1eA65tRObiPrI192hs
47LkdW3R+idhNo5NCD9wJF1EowE3bEEyJ2KUTVY3oqw+8LaTd8sTqNPWaZ/3
yMm8CgC08rJ1d6tt+eVxGDDGIJDiA2nBx8HfQSd/HZLna0CRUvXg52DBPiwz
YYJr2pAkeq3FlRPTuzptJNM/99MQ8X2fo6VQx21i2yTKwTGdse4t6QUs6Mh/
Ohesrs8feRwZYTp5vrLHNAvogW9vFDVBIx1MYQZFq8MN9sA5GyHNrr5knCKE
hJxod6h8Yb1hW8d027xSrICDCFRmfb9wKneteKxaBR2Z7Sg4MtwZkeV57DjL
16+h+v2pCn4vnV+7dQGgfQe8KwREieTkyofIXqlGYY+t7A+8FFUdIdmw1vfi
HcIVXYxRN3gQ658ZPmiIaTBUa7PW/BlkNBkQ0aCdjXPHQw3tizTjuPqhPk2c
dVzFMl/v2OPN+NEdKvDzc0YfKGoiLpjgHaTdrAGIxVX8QwYpJe4E3vxiOvwJ
y9e7MAamOYDHWRE1vhoMgsJFDeebtxmaQpgi9yF5LXciIYbLAudU0Irg/znp
ZXYhFJldLGOJ54HXghmUth/MCcCrIp4P2179A98SuGmer5SKjC0OkOrkJcQ9
aZ4CukueqWR8asA8735XVq7/QOyA9TZU44LxGrNBaUuMffL2TFLcRgci+AQM
9moQ6WjCQWcqdibrwZ86gbNuG7/Yif19VOewTyYHyGm+DHFAlTOeRLgXwUNh
J5ed8VSNEzT4AzG2cZavjuzAtMjuhKq1h0+Xm6d7G4Repvs+AwRDiZt9OyUO
Tf4Ibxn0EjcZBP76q8+t6dNC6KnHu4xTwoVQnExQGVR009fvDSHxT9oEAeT/
khlBisrk/mVwUZRIWqggbh27O1McxAtgOkbCSPUjsovva787dfUXzVsdwGKU
SJrWHjzC5OP+vyoBRQ2tbneXtYZtyFoMXIwgL055020rKtCmIKeupvEeBS/4
uNCITezZD6sAzNagq8AkM/Kv1x5+GVjGKzMf/OeuaYC7ULsx8rcOOvY7GCma
qNzRkmIS3oJmuxrfkckKUOFSlyIklhIY5sCYGpXMBOHM55Vexf4QgfOPRoUp
VtPeaq0rCGnoinbE9pDr7a41OEpmVTlYn76mfKhwZctnUqoqwdY3nEahbbmd
0opxZJOkh3mcHu8Lkf2lSmm386sZmWzmsPqVK+zihO3sB4A3wf3gn4HbvmC8
HPG1SdsvMUMJfTxQKsD+Ve30xDbz9pL5rLnOcjjWo1dbnUwWg0NRkFnIc9LR
LqsttQp61v3pC7E5GPjMOvONFrSqFTPWWonAAHUjTKc3+Inlc4uCqGZvpC/V
00u6RZqYq/BnPR36F8fBAzOxbKvHv7AYyt1qkuroPJMX4T1X9+kRurSJDU6S
ZmIEDc1A3TwRcjds7VnDjgSfa6tBvHLbnuUjU2KSjwWCLdRNEKFxudfaYwA9
+tEyZWsU0d5hOraz2q/dQjfkT5XMS4YWjAWYOjCbQaU8+z5hQjc2RQoxa6kf
2L5htyqDL2mQLk5DKTQ8mnttRQuMO6ZViWJdq3QvYL+D4Xl0oeCgeA2XcscX
bAdUYTX5FnXFNerW58MrgxWr17QU2pmuyx6mXB/7GoZrVnK3nAZKxhAf3Te7
ziQL9lhtwibW+0ZO4F+WtWBehyA9AzHexf1+Ue6sBISfnpPaaCtj8He5C+rS
vS0Iymc21llA+twkD1WnHwBGyouYduU9Mm+re1wSoKbufip8V/F3GlxvjoR+
4OxVjhRUDqPZ3hun80C8i+JWsZ/T855+ZCH+uxHpLjmLTvZGEeVAaYNK8J6O
Nk0mc8jwWdoe3QzsvE5oLRaT9AohP2bpVNJd068LI4Q3i6B5U5v7YRv5K5zJ
IGDs0EkSasdCc+Z4SqXNduPQjzeneRhXtGWDG5SZkhIPLvb7E3CfRMvJBr42
XlMOvYEuoLWYGbAqZZ+8sHWNEYVgTx/qoXgv8bpqI1lFSy8JvwWDoQsqNoAq
x4gnyLssgTfohIAwK/9m68/bWI/aOgszxEeMUmwyfFyNeJXaTqAQi7KO3tYH
TZka1iZcAUvpzGT2dHPOZ5eHgPbHh3vdmxDBiXM6pz8F1XgPloL1337j3PaC
RldXbyIVRS7frwQJ1oy2OcZXqj0kXtMf/bX1+EZ0QCUKBRV33MY9xZbss5AG
IVHN4H7y22RqpfQoE7l1fAc4QNfIqWdeZPjRqNJDD0kpOhm7Y2VjLT1uBIpS
XBTNUZ5roHesPImxdVuFoAj8+jnjw6HU44Yl5kCZBtoavr2okmxccOPZxtZW
H6qLa2YeI+IF3qwnmqNHRTxb+MRqDv3lbz5u5zYotuOe48Rm2Xh+KnZHz95/
Q6Wk6g0wyFizeTgXkcgb/2DBexDR0YVFFrc2OcRWRWx8ofW89uYjxQzBX4i2
1o9evLBC8c4oQXrjFEfbToKptRwFzX/4i+kpt2KHJgFkN+ZWBkh9dHcBb6lw
4AHsCxfI09gzaJvI+Fdad8Th5FF8ReOtMYtVQcEOzADnkY60FXzIYPdr4qur
uBzZXHDb7j95yidLlGT20NhNX1iKj6AEFr41lvjawGRs+eYE338gYnG4goKA
R1TU1SVk8kbzM+NkI8tj6zNm+GNbt8IVFCfIr1xL1vOFAikQ8S53xaSolOfm
QJOVcefUsCeBR2FIfnB2inRO5vV4q0P5q2qxTHsiwlJryb1XBAMXsq9qc97b
Qgg9vuOilpV9HieuIfWPRraSFZZPNvZssS4jmbPvq56pMW7twfyhgt4N6tfT
GBQERSuOeNGQmj654W0GzD9tPQcQpv7dIJlXKFiJTIG1Bvh5C9DKdQavJt9V
mQd7qYmPEogqe8ycNzUT6EOtOvkFBDnvj5l2kX1HAvmWwOTDG/0BdVtcsStp
FRHynpRxXNM/1vV+4HL93yHHhTt81gI192newZWsTPXOBMnPO95EaKXxYPBx
QCk5+iGKYlYRerDSYmENO8sFXjjTRkV9yhf9ISJrR7hcsZjtzX57rFRxxXAE
Ke1zviitimbAdkqjBPkHcMpmFE7B01b9VWJJ7/14zt/p6gMNHmWT9vixpBzf
ucM6Lxtq2WCxcugWekEWQZwh5Muk/70lgpe0R86t1HIf3Nhk3xMPPebwlzHT
7csj+mTCixH3pMcyOFkd5V+rWeCUhWEgkUQy2kk4V0MChQtMMwNRtkORthKo
MsRvzBFbC1RfYEWKc+a9E6jLN9C0OBei8M+U/VeUKj5xPB/RBm7lkXjWhhK8
ZZL1Bo0bAQpdqt/ukpeo0tKwrr3LxNj4HTNSDVNaHK36BWcmz+fiKhNLDm1J
XUtIhTlgqOePdrtkP9fA7ak3qhBTjUVu0lEVSv8ox9RZfChOLNGOJZTpa6M8
epJ8UisJMqbkEOw7cnJZMzWe8Kzq+Jzwmb1w9qPdrV5iWsFYI3zNvOm8DXNs
xPArFsRVZ2Oa2hNHs7u6byQ4Z5+lZCHD3H2ultDQDkt7VhArHrDp/WB5s05A
STm0D+sbTut89sJWrnHGonWud3phSSqEgPDBlf5VL9187eYihzI8ToPCGoCX
F4+3VYdKdTaI/prNvp7g1l9BuNUBAtTPoUt9QDOhiEhn9g8ZqdOmEUvbjcuE
ye2LKhvm1bfgEQ7W3CfKpil5HJYu8sZmKvKkgihc5KH/k3nZNjSBOjklode3
4qXk0SLqahdzCdfHiDWaF0h0VGYPla72mGs5Va09Dulf1SPlV+gCCV8KX6lY
BQNGhspYjHm2LFilQX9IB9Y4PUZOJQHPyQexx7VWYZV0v2/REH8VvxtSnuDa
IME3LirSKZ7EX+AnnGbgv0I2KXRjyomNNTeohOg1bEMKbT5nRJc8I58aCpS/
nHhBDoQVO/YRlizfez+oEq97HZ/t0GLCk3kaALTS6Iiz+71cdh09nhxaJUcJ
lQhqd5jNAkq9i9Rw/6qQ+cowRw8ZUcK6GEtwOeYlhgvaATW2uIjabpS8YU4b
KAwdWH2SjiscGOlaRD2+g3e3EhWiu3XaembOERV2W8wt7SrDCOvPLNsY2fO8
AZ8Vtnie1kY1H139CkuhfBWT2vDENi2/GwNr9ZZpFdx75oYCziDZiERCVUzn
huHURVk5zm9K1YuKDpEqPPSU4a0fu1S/LGptD0c9LfQYMJ6PS5On6g4CIkB9
uvGeDeDk5xXQ1yyVtGHwA0Qn6gK0UC6DWdWXzlwLH221TOwZN4HbfsPpe8Nx
ToLleAosB9dJ2Z8DC+w6YW9HPe+TyG8rXv48XoHi2OapeAB2O98uzZ1otjxY
NyvBcI7L1x4GupvultFsTWYzFIcuyyXMU0926uKhT/OoodzRwFDXQi5vlbit
mq6QYWUBjwIkv236goC05Yetuj/cthudBAlN8k/6l8Ft3dG060rBfTfkhEeD
hy/b5V3DQjPASZ0PJT2yX6jGTY+OioqKaPegZ8jeVrgsF/JcdyMdbyMGOb0c
VK0XUXM71ybDZcw9/mJ2C83Cy+PO2MrDiX7kyKJ54Y2F6fJrmJsSnCSiyym+
LBHPpdpIpirxaFgo1mK/Zj+iI9o1J5RzP1j1k26YYQIDiwsQpj9qRVcMaMEN
ErhQZZK+/Fr3FpUk7fy+5tyKQSfd3Zh4cThBjAjohMljb7dAv3qZw1+cpf+P
EU3WJtMvc5/vthEWbgQd28dK9aCbwT1C19sQ/am4nbzG+E+6P5DwqXsHI9d7
EsiUKGhLoLtP6O1S8kivyFzupKLy5NCNxfl7WFDracfjsTdpyXLR4Yzq8rtg
CRrU5NJwcNq57rPJQ5i4EOjuWj9aulAT48Lja6XfySqh0ppRNf+GkUP0vMrD
n5c3QsZhhDMute+VEN0OlHZ8h+O4zGjQdKyWYrf71Oc/O4TaqJeNvdh3nVad
3haUjEUHB5iCQXo+iiPWUkcHkObBD4aA6F6gvQOfqRSNAz28mBb3KpMBzZST
2ye+6nfu/mdHEar1/GIJ3zroRb3tugfvTBn53vxWZ0vPXKfVFYhYlJAkYIhS
pg+DnZuBwdb8ZnuSc9QawjHPdUtzaVo7nmih1KGAU8z/Erq6FqXVQn++YKFS
m6Ev3zVQhSmgmp2uyNElf+mkPoKUVT0uLkKjDrDtiJfHbythukMm2difSJ0K
lIkOOPuYzkYKLxxBdB2vVhcllYVQ/PYHVFAR4RCyJ/GbB8QMbZs5+yfNU4YJ
LbDb4YMIKVh9ft5id5/Ph+IxXsgzNP/VB1uWKk8ZWOeKTD0V74rrDLGT0DK/
CPrGAwjcj4afdsVL3ZCDRngFacwhtE+ndGYhMNp5RI2BE0tmlzq9jMVrj7SC
tw7XuKaYsJr6JZ30dG2QLPjYePs5x2EOQuSAD/1cMLncBxRlo9ND6fTMXJNi
O8hT8f3+NNoz/ZsYuKWT6Vq3UGSADyOrQFjWTflXu5X/yfqh9xEvcw3kO6QC
qneoc6iw6s7XPBbZ1e2sOvsutLSY69t6c3MixkDnV60rKKhFIP7H2jQmDCvD
9fETv15+N32w55XMCLMvyN+KnWb3JaT7AS1sBxe5Ww/f7quxt0yZcgbpzB+k
XEU13BY23aIDmMVkJ75nXL2vjRejNUSxuTMqHwvjOahCKXnmT9yIThkU+PKR
4RRx+Xknv/rPWSMoutqVN4c7dPU6ynBiUl726QI9i4SvGGGIpEwMALeu4BeE
CD5wy803AgMV1gdlH2TEjxEuHdxq3LCL0ENYc8MbGMSDWuphThkPbUlWGlpT
kjn1X7tWcarGnOVFn//1Aq7ccHOyPVJ0dPEHLILOTyxDuPrOaOc6xrYXALSH
g3PPKD4mxvSrZILVWkkl+DPF5EqkUgOV4cbjYxukkbleLzN4UpqwOlA8CyuF
iYwx5M74IWP1BEpwBeLefYGy2MSm942hAf1NLy/bGmRem9cJ9mN/M7qWLIdZ
WFHaC97w7UiAKGHZ2OzpYCGUZlh69MaADugc3aDsxQQTGeVG3GMPpguQrhlV
e8WC5j7crbrKUWAa4CMyb1cSiUI4XFc4ENcnVjvgamSrY9Oulla2M3fGp92/
WFp+Y6PL96eXjHhd8wIZgC/O9IVEYlnLlRMOsDalnKTx4Na0HZ9PnfyAb1Vo
iwkdSqRZwKQe53KTGFGhRTVKTnhcE2norRyRgYx2nrJdAsVh4ClWq8NbYKNu
6srPW7FCeV5wsTSRB7R9lHO+DW+2WV9f6u5lW2C7hVc+Tcl0lpt+Ccte1huT
qtscmdxvHmfbO1cB9p/ru5vbcc38WenLbb0DfLwMzWCdvtaST/cGr1IJhMyg
LtXSCvYnp2WUkVArg2Ir/gRujL5u0LZ8cj51uz9bMS+4fiBNvEgUJ6jVQU/K
WmUTy6NaZbYGPjLSyfk+/TcBMPME0I3Tcdc2OkWm/yDs/rjH6CgelduQ8JVu
XmtrUTFwAMQEYa2DPPQm9Pmk2OOT8TG7DYgqYXDQ+2C7khotb7KXaDRkyo5b
JE5PUd8dqTN/MqgYpg1e0IHTQo/Dstk+UtAeETQSO+73N38dhlBn/vJ+URPc
NR6mndDz10cVM2/IzgOm7NLjwG8WbyBX2NVrQxyUZT4oHLcuw97z0jvFvmaa
5AhuLX1VuDg6RpzF/jBn3qzK9Lrr17AiwvIsIQkOfiYuXzg0G92fWBjv1z5e
HqAPhfRsWh7nnryi0V4jGb3Kqwk8tGEncAGZO9sAui7XlVkBEaRlZ+etAtyQ
v7fP6kc8Mu3iMvHk/YLY/IgojSDZM5PBqR9Z4mBG4AiWARFk6qiXpXjFK9Is
tOkdcB/Fae/lDya6f2VJCGTL7ZGfBOQkDjAnh6AZnunWMwNHK6dj3hE6Co71
C4ufuNBmadn9W+djdcg2b16ypkD1UkMV2YzdRP+aEalHuH0pdbu/Hfxd33//
U+Tlr0dNYm1lrxj7nTHuHP9ygI+hbsw/V3vyouppVGHTD5KFZ/rPjXoMpCEy
Kxn2E5bvfQGo4bzUDMhlFiKUkv0YfanbeVT0pM/ichsSG0YbpEEwYdi9PLqW
BTIXTrDn32jOcFYB4X0p6TmeJ5L9OPR0ZeQqNTdots+99pULBBpQULEqc5p6
+H98knuYIT3UipbHM0MlNcbiYS0bWEx3EaDEziuIpBt9FkIMGB9VWzqndFV+
QOU5E54KubQ3taSzVKWCb6XGI46sFJGRer8fNaakw0hhU1tmSaetcgAXP9BS
bt1qdhU8CJ7ONQtsq1EP/F2FYlmDX1tXKnaZmhBMBY3t3p5Dbc5c0zOQQ19j
syGR2BO4gC8osTS9YfY//hqVecXXTyGlVA/CAyWbva7Ws56Z8yEqnMs/59uM
/DHyzU6w1Yqnh2R6HJ1K7czjT47HVymyJYerwt53wexOK4DLIboefIfsYRh8
C3zUsM0/Kr9fBStHHSwpqW4406OI1R0OLayQ/1/nDubPCiIusi2bg024JBgz
3V7MSzpCz/HdsrysE2Eul4DLlJSdyww0tl8vd7P1itLAsg/T9mW5zSfpLc3R
6SbpmxU+G1DjAmF9uJWwjOcFaHFlfgRsT/ss9YMTAAxSed2HlhW8IISnM0eR
ExI4q/anr5U0vmHvLifvVccfpYe/G9bMg4O/mRA85wEEXXB1B3ywVf7RBs5J
DHqO+4LiUrHysUJEVENAGyaWelSY9kksTxDeBI+sjumHG5EkkHo8/w0f0dyT
yHl8BPbZnjBcvDRigtLa7timacSfFNQxcutLFiQeIBHO2XY1PJO/8t1BjxQF
iF8BxHKlzc5sXqjtesrCxbe05DnpZUCkwQEjyVLReaoEQd1sDyi+rs+Sj/Rw
Hovw2qEPsjKr3LvP4n02JQJ2qdSuTOckjBuHpEP4EqcR+fwobvoSmpEcgvNA
3WD1b++XGmHibIlCP4zq4LWd9Up16/+GsH8mz1TVr+V3l7m1Px/AgwO8UkhY
Ntr4Tc/G7stugc3+OI7vWXsuWdZdGEUbVAANSskW728PXJSp9lQV7hDY1Kx3
he6fqgJmyokD8FKYOOcaOUgEYAdHmyXqsCaEKP1N5DyYErbudnN6r+o19wE7
DWOdaQKsKNhwmuaSZ8BbNSauDU+t/Sqslw+URSkAbRxqcHdc2MX91dlAkkFj
P2TUwS1snmktyf/sSmBKeM8l5mF2E6nJge7ywLTPnluMUWxU5vAKcVuRn/iw
qlCfJ50ttSXaq0stVZdejIedx4NoN2NOknFj/hmu7fiiMTGSh25yJi8F5rli
yE6L1+sHJ/FVA2XR2OYj8Ws27uk/7tWVHxLJywzFiYpAcoz5gSkXp1oeCnzm
LIHxtOHZzI1jyHG7g4mXQaJrOMcC9wlh4gYpz7PyfZgPuaxQNignVXAtEkxB
g7va9+0PUFXmjHh91/1xhubSZGWB3LujY1+SjtS9OYNpbfFIQLkWC/9zyQ2v
stcFsX9DlisJfEc6/OlHJgKI1YFqkGXe6x66QOpNkCVowUxhkYgp7bxkYubR
00EvNqR6qfRS+gFKMZm/AybaUDkxHtSKbtC4U2p4Dh7JlrylyHFwW5F3oHQo
Meb9tuDJFeXD6GAGGATHgsGsoOt4kdGDH3rtftdFeAZvibh9SZ6jGWLh9al7
M78hbwzFIoL7CkMKVfihUO6AJdjaaeusJsLKV83NSTWwZSgyrLN3ed+EcEJr
Dy948lNNc2+u0D1ZtwJaeriToxrqUNOhaTepe8Ee8pcE4zS/7QY4Z6bWw6DE
x+07rCgiL4NWCkt4xuUmirfeIh+SDlhSlwghGBYs3jgPyWuZ3FLbiSP6QLKu
xol3GJVrwa3hWU6EB2qpzBMdNoMpsGytyBMB6L7Xz61iZ1EgKTZ3LCVZh0CE
u5fwCuPD5Q2fOACj2KvVDwaXMppUihg4sld4omT1gyTBEnKaLJXjxv7kHpjZ
a+nYlvwtblnz89hhdiF8kC9HE7BuflyaNMzGG0FaOONOfx139g8Dson3WkBw
IBlnkoPZBQYurFBuSlrIRUL53xZXh/pScbiKiYNe9+2cxDAh+Umx/rYBjy/v
6WA8nEUhW8Ol0BtdbGmR0KUY4/4afMdbQ/Q419jxDL40tY6lJfGR/TvV6fJt
2hn4GANJ1RFztr3EV8zN4IzmzElFVsVo9RZ/UQD9p6WtarkS6GoKQhyvzSry
KraRhrFgLFL5YrfLmzSZM/2MwmQH9MoZ+PtFplHS28RrS1mWzWDFK8qLpG+i
IYk7OjAgbi2BtEISwIoRVRqlZmfBrijO5H94AQf/NagTReRE9peNtXc25AKd
biwMM/wck8pTITH0MJ8BOzGsIjhPGnZCH/tsjCy6IboGvzlN4gH/QzJSrpjh
8xoFy7R317U9Sl6GrDOlh7Wb2KzF794mAvvw1X44G28Y+46oMBp1D47Y3+sZ
/g5XetdAJAwCux9GSX0C7Z7fWrXJlvI5eyV9id77Z4Enke3HoZNX5/B6dB69
pOvIYPK/h7+VBDmSXA8tbESoEf5YfVqNFR8Hcns1hj6OX8P8RmT0G68UP5XN
Q9a7TtGACH8O10isX4EUeqGSAo0zkGR/NvoLfFLPH+nAbNpGKMUvMIXFDUlA
VmT2HnWnRc51NJ6H7mO89KLMADqRZhntG5dJkC9XSeeqNQMXwHfqlsb8wxDH
7F8TZ3lJRHv17Rf04ccyto4Of03wyy+kWMoNTdeyjyXi+W4mk138SBRoaHY4
DDeHzlGeljTd2MbGOBD/OmSkZ5aBuSiSoWmnQl1cDROnbB2aSb0MkbpMefoy
SeUW9zoV51Vb2TitGhq//aaqtrBrALiDYFY5DD7EoNSHkLrUvGZGH1QElpS9
QsERLGlScDr05PgooEAtq9MGy7qyW/5dAy+d7h45mHvwMfUC9lXwWbSzi2H9
Vt/Btm4EmTSfCQMcCf13fpd55uyJ4BSD/FDD4sZKuieANvVxWGB65tLIzUNw
lpirQuKuRVdMxIbZ0s4jhOOrUEchBh+3MzfzW1FYZGJVj/TxxIcPdMSiFeyY
f9KkIlDPmt8bkex9jz6E4Pjj99fZXb7sckd4ydgjRbzvBETfNIpoSQR6YMnw
1cG3KEw6H+4UKHY5wtAWHvDFWrTdlZmvYiWy+XPHe0Vg8DC3WHHQk4xIYu4C
DwwOLn2236USXLejJmUGZtpLGM35hMcT5deW9eTSSSaqKvFQ3WsveG2ptxAw
scaW8/KoLUfgH7gLZslfcreulE+nuJ3mrE9rXqHbKfyLL3PyVeUDH1+v4rvU
RJDi7SoccwpEO2uC6zpg6WNzczyzrqqTNMwz5svYWWxyH859tkanje3qj8CO
O/wqOVbFTIJRN0IasWx5OvKWLPFZXpIAz8JcgGtTdLn0m63GqhBGCFuHQxF+
DHiQ2T3e9k11mVaeEL29w3s8+0M/9jmhOEUSHh4RXflA8bCNbIILdhQcTaYM
DxjdYbVU3rkV7s2IlW7bE38PiLzEqSBncq97wPCmr8KeJTRTvdyi/8X3XGNS
mZYR3/kRv2V/m8U6FK9lgVJZxWHUFuoyXBn+BfFItiZBnYPEu7JSfEJ1zhFJ
wH5I1oycovNNpk0Fxvpk1lWH6wQqcFAXuMQ41di+OAfZ2AxXxwx9O/WxzGVK
ebtTm7Wl5aj75wwkpbAYbtA0Ms3D7xjtBqNqO0JhNtM3rTGw9nel4rKk8CiU
20jhMkcjDILRVC4adMKhZwtb0HGr3XD7Ois0sFp6NoM6vZUqZDzKT6mxRdW2
8jgQbvNLVMcQLbAtK4zRrnreniSfginWccd0mRaXmYZ5sN4bcTb+68qAt1Go
Cl+xKg6V70/dyB5PCGCRZ0aLdZubwsjiaCmMi1vuUtynF/2Vf++cYc6h3nup
fN5QWWxHjQzkfkKhWiDaMRuO1ABhvMoIPf9AZOdKrOtDeLpwbptF4tXBOg4d
zmF2cFwGBloVtuN8CZZXEwgdC6V7GJ0iy2EkYO9JNnjVnKfYaiIBWg7x2UFb
wByM/BRo1oxBD18VaTQcYl3REwC/wIKltid9oQwo30Jju+XJ3QgKuRGQpgQL
cIFil81+WBpyc3VaRIRW4nPM5veeVE8RpMHsRElcRLvBN5eFKKY9Ca4G5eEI
4X1XW4XAgrWI+s4Goripsp7vC4/oKVHs5zaTHqhevb6ytfUHRhAqXZx+uzlz
m//9OOBW8cGzOCBtSFpcQyR+hxK9muRuHk5mMhwwIVwP3kIhO8wkacMS5J0v
etQN12iAyA3NydevWfoGT9WMeivZKiuWrkB4NpHiaUkge1DTlGL0MeGI5FT9
MX2TfQ4kyxfmJAGxlp3DYWdqUW6qG07jRvZXOGmJhNAsNA0LsmRVu8F5mJGd
ppIiMD7SPxgxVFyPWo2aBWWaHQzMnOwKP47s6qIf7PigL4AXTutRpydlcLRE
0iZt6Ny2saAHaggIKrFAHoSvYa0WK+xSwaYub88e8QVNp+5ykF8dVf7pPzzk
HxFv6A+/pqL0eBv+jnqbF6kyVLDAKOkg0fi8k0mlB2hT2nYOi2DviCZ0jWqh
yhT9bluqj/4uVI+vOg6LmOYRZZMNO1jseEr0LusJIW7UrA2WDKUbw2kLLqf8
DiLYfDXgvion3CyBHvAijk9HZidw+3qZyh+8i+AnU9KjxymqZ8jV6ryBA4mJ
PD1ZiaeIEUXWIspsjIlAXF+pDMiPeGNuBQ6Q8mVvYjNzMYXitIF9xF7SbAsG
1KDEijIJVY85vlw+gJEkUMjlj3WzNEAHiTYz0ZlFxqzHs/JFmB3DiyFS70to
SGkwOlwx+g7yw5tAh6Y3e7Xs3IwmIa6FsvfJdRKoTmT4Px7TNK8I5I/R5vlV
3S20LQrQ736EgjaPT+a8dXVK/BzGXn9hDRoEUFM7+1Ve07NrgrePDh7pwiRE
s3FThI9etKnCrwGuK2M4k3ebyNS5v38YRhEDnbWTd94l+k4vecVxRYRfqnWk
9K1cloQaJzXE68xTORuJdMYRS5Ubm5y3gHoE3dUIFhuHsKJsmc6TKGQo+DFN
8FZryOzV1xYydEzerYkdAy2xafLp7SS29smBrXa3MG68Ki43hmvnkAbtGJWT
VDqeq1mnXL2MkZwqCyAlrV2SZgWaNLCHKUTNjw/gn7h3Y5DmNOA92HpNRKq7
HGEC4PCFXHKFREIMPMf6Oem5Q46+TxEIPaHZRio9VlW4XLHU8nxNMpm94jLf
s3Cqfw+tamaFjniltesUFmWc7R6qs7JHt8/JmHOPQsW2+9fgs/rIMPEL90wr
aMGJK61is9LirLEtAFysViUXdEkn+JN57nFpFUCNEcWsq+tHvROyhYg/cSeb
25THTcF+M7qEJv2z9Wm+jXMLJMGk39VgVZdNTDNXc/4m+dL/0FnKfPH3ELhc
TkAtt2F/HiNI3J4hIFrW5EgGc11IEbjytpIKEydr09oeA0KvbT2dpG5zZM5K
MGrhvx/nJHiJkwQcmvUnht4aOwV/fDU58mncZD7+ui0L5x7nHHDBls3aSMra
n1tgDHdz/WCGcXS3Nbb9quV1S2SmXXQbk6V9ZheLATRK32hOMfxWnYEAGR/0
Z0qIJ3LDWS3NHWEbVrRNm/WG4UspB/T5uTL4mxxAeULJSx9TRPvYsgeoLQLt
WLmuCnCOtNhYHLlqYfLCZQcblhDvi/aWIarHSaH0IkHFN0R0IOBIau6Dn1DU
LbofOpdHGlBOob/1IrbcaPbTHFlJA4kIdziBmV4nBI4GkVXeKa1gUcXs9IM/
L/efV/WzPf5JcB9Hs2PXcFL0sUHXgzgF/93EJzXWTS+1sEGTymO5TLK2IOS4
obtKdQsoQVJK4gdrJP0w2YvMT9dpW/pJkhP4SRy8YAa3gd2x1QbJSTmNbsA9
aedbxNSn0USOkhsqLjYZJqrdtuIOkZkDL9O9KcxTnHQa5O2dbAMb2mbYFxDZ
o5lw7T9LmGqpb8LeCt7HoFe22XkJHT9TuiLFR2ne43aZDO/8ijW+jnlR9Wj3
Y/PjpUCL4RM+crPFgUMnDcDaPXqKM7gB1Hgt68u8Oa1FHdFT0BR2qDCQLgGH
ZuO4Rg+NPoDQggamIuQfVAKaCbqmAznmbhX0V96xodPd87DGd7xM3srs+4Rh
xM848+hQEDh8ovoQcm/yjYzDSPkDvIHqzaDgR3oVNCUwyk+t2Mn3P+7T30fs
0BuXsHe+iv8noIN8PSjdWLkxm9j2ltRMWtcvF2o6FNkU+3q7fhJ4iQne+Tik
LVDG3PutpQ9sLlb2JCwYWnzi31nBtLr2vJ7vsN9i3Ap0PWAOe5qI1S9iP59p
RImVGssIO7f3BVkYo30oUNYjByk5Sn+F4gTOjLmldxq6TsU8R6nB3v1X/QLC
g4eXhAtx/XNcjDs1x+y4Yt4xpo3mUKZ66mAf9bM8vO7VVfHuuGft/vYRFFzU
1MuuB2ktlSmBuI9kmldutWCxA5VuS2CifpDH4kZi+xml9tAfPKB8klxnvC4V
LrlLmmme6sk0VQU0vmtgPROlOeTnutPVknIjISmiy4EGlenizyjnutINocUG
Ck7qoNKktAe8t2ghAXaUzk2d1zAMlYbz9jZ/9LlvDvXz5Z7AD6MIQuz5oyH9
qfgsNXccq2kdyPnFaNLZhSwyXYmhcM19QOlb1fOy6qEw5b0fYD9xIBBcxY+n
GTotFloR/vJxFof/yPV9nH19cioZ6KNfBb/0m5VLIRQIhBQxK6426JHOzFsg
fkhmz9uFZ3XMOUD6YCdipAbwtLgq29WPEpElcro1I9mSGmi9PmKecGhl4y4N
UQjV538j8z+kmr2fFVI59EWQbAUhvJ8g0ctb7s414W5IvP28bMJ03avVjd/I
7EjIil1an/orOu35pOUcdNVKGr3MB/IOVYB5bS6lgFCys+HeBR2pmcdLUHa1
k4/p62RU/ThiLaXf6s87jnXRxxMnf4xrqal6Nk8W+pUVsCfgKz3ymQYD1p8n
E6FKumqzLd3MXmgVRq3c28yAXpL02aa3XpaK++2ocpp7XTXNu+5E0L4VUYdq
Z8vVrxv5JgiUzcHNDR7j/WsJKvalMrMCSg9uJwjLi0yufQz7ehjwT9zPIxNN
3gNJVpx2OVVQlnjvGfWwvagDs9bkXO/cpuJYM2bAVKvghJumXSy2fnsRsLvF
w4hoqO9hE0xTkeCO4xtVyfx3DrgX+bVwUbOf/ggrWB8i9Mgbc4ZsvQ/w/WW4
ptzWTQn8s9Tauk5zVN7B8Slqc8qkZ6++6vB+9NOJoP3ajuQCAT7Nj9C7KAhj
daC+q9zWNSSotyDQYvF+UL/y97Qxi+nE+Kfgx72AY2WiAKn9ps0AcoaovLWr
DmIavNmCz+GK30dQH8iK4q2yFyJ676j5rooqFEW6LA2qoOrJpu9m2fzvI8gt
iU+o6Tv4rjMrvgJb2VXEOKk0Fo+FOCzMA8HuIM9/+B/ayI7/+ov0IfrUdaoy
CvRW3SNLJL5CMD7r4QL7CYyw2h6Ltx3Tu5hMiZ2TsdiCicfoGtxoV1MXGuo4
7pwWFZOkK1vSgzrNNUHerj9EnW5eEgugw7SWQUoO6KT1LQB/8wEwsdxli6nq
3DUrcG0I469Aw6UKWHA7tGUL4IrRfZ9PnGCoyN6Qej5syjmtr14qst4+U18p
xYkEbh/639NtHAXBy/li3wx73g0EPYc1tF+erdCbFhwavbePHtd+644bjbE+
y9RzWWp6PSXsUQN+jwpF3CcTUeIUVeWLTCI2gmFX7PzYQ9qUaBUL1GAqW+zM
hX9jEoekiMMWNAd2B5tKgrSh+hUCAtqSpATQAfHLlPCqcSUqCGeLeET5VG9+
XK0QBN4p03d09Q3YxZYQ7QN/RMJ53IITjNgbcdg8Vmayv/kXvSuPsYl8deS1
mvemp5F+LbBiZYq3XEiBeBskkJ+fQN77DZFyHWXZPujQrc7RoqiLBMUHEynT
YU+nODowv2HURBhKTIDhDQL5bTKVIM5UHNBYWdMizH3LiLKIzgcxRGfLJKd4
gqsJ6WLqOM5whziZpxkxe6XeopS3gdKQR46MS1Mf0xbxKck4NZIj1WhECAHJ
r8K6LATeikk6Jj+PKQU0ND2cHDKFG1EG8xbG0IQdaU3fePtpvc7yq7O1Mrww
BfnNoTtqJXYfADIiQy4qMNDjMALKqGHp1t9uEvaCRmKUL1+LZdVY+BwpDf7v
7ojA7S+eFBPo86kOaFvRr1cwkSZ1j25KuUm97a7NTg/6F9mGrfmyL7xybeFj
LXiVS3YSmMGBpaWa9ffFdNUHlCIusuIMLei8mmkxEpT1RcS8gabKksbO6CUF
EyQZcc6zkkFSxxwqjgY6Y3EJTSinfdejgm8NR5vmqB6fq6+KtOLMH6mzoXKt
SfI1/unaLsqMWu9Y9TOIO1PRxh0ukG7H+vvDgf/gDt08oqiYgfwcZM1Vl56h
difBInHCbL70ddbu2LiUQTI+ex1xT+vvMG8ldhC7Z917Z4nfGjB54h5j+5dy
3WmIJ4BmsDZXRsHmV0hB5roy39fI/J3n4rEoz73/QtCPdFrhDZjLdt78Jgbe
lQMDLgV/HisN7aSiWdAKHF10ustxFkqreDo84hXqMaUeYuHTsshnJFi2g10W
O9h8HJ6ivoFuoENwjInkcA5o1vYipPiyaws/sPs7uBjGkbQ3yc1S4JTccKUG
e9nf1NiWGanTLuGLkmocaLdmAbNNkKhWrTTx7stjUf6rCbDbwZe1IQIBXd2z
64t7BAkihgbZELKSnbIk2Aq3V6/VBxKo35ZNimDhK03+5eRG3smkPEdqVe38
/8ga7rTaTa63FljbGuK/y2mXCw2CNA05yT2m6COKb9T1n+ewGexpcOWvHrCX
yISjg9YkOldi3Ju24Jid8pZIeQ4zMn2r85o9CR9j8VIRrLbq00OvsN86KOy9
C+cqqIi0FkIW15imugZtrVQmwdAy0aEfws8LxazjBF7cSo7ZIAIG30L6ncIp
Ful67PE3YMqQG0RzgYG+v0HpPJDTQ/KlhxFDGOvdIn+BP+fLdhq/fj+EUt6O
tS07gFmxhx6SNGXJi6NXOP+F64SiDV7Ja42Tl+k6b+2/UVcqTPDRw+UOP4d5
AF+1HgaHMXzPogl0A/+0WZ4jR11ViXT3yHLlSSmaYBtDK+p72n3P7iY1vEPN
t2TVHjsjmwiSMWIG62Ii8XNXJWkrTj+JxDt0P6RwuNtbtbiJjtAqnmAbLKIX
fgPnDnYZDtSoyXFhdW55F7Wo97sLAyjIoG8JMpyswPCxjIoj9Kd9FS9ByoNL
3R8UjK2XFAyusiIGxEQf7hF6WPnXAFXl6hR5IPqTx2phzNX7DV8o93y+cNhh
geMr4A6KpVsGbhc0i5u4XcOB8il/uhVi2LuJdlzNHfkOb349rohnS8PiiL7E
OK88JUBdaKTKM87NiLnTIhv0hem9IJphvHAa5FaH2OCDiCEbzw6A5Vp3/SDt
kaKmNtDYf1nVdJ6+rmspTTsc5iXj1511Jl0U8mStbVRrgOzWZkJ/7fd6R4Wx
EmTLGXKKuuRH0eBlLBYreebrxgIZaoh1XzP0ll4AMTsnc05n0HY4W+6jkbJw
Oqbv9Kf4e3x5CMB0fZNDLMok1trOoefJyPVOpAjHAcwEny+M4sQH9+dQAag6
hCBKdU+w1+enzKBdRMFgEqEimeEh5P0fkGFmpoB33ALXvOOEbsI+E75yci9F
T0yWXcXdwikZnVl1RbaUF3PFR3TuQxer8+j6Ygf+2s1F9uO+wV6o7DGP7412
LN888EOgX4/wQ1HA8hjRrIfMsFwy8Zelgf25OOd/R1b/e5mVi7vRDeTuR51N
YhWglAdRWx8H8cXyCx+tpWLtFE6U8YyDGjC44KXYD32wOKMzWyUX0AwYzgaR
jiPhdsWdFi5P3smqJSgnczDYzxYD1goppPzfATbUJ1TI4Zya8RXIR2QfA+f6
hVHS5yvfJs0IAqTnfwjn+hZfCPMxA1hDH65A15Jk6K00jaCZevuqfjWMk1lU
9Nk7OUkC+hJ5tloVI8S9KzSngHNpRxaqZEFCxwIECz83Gz7N4A840m17N4Gs
qYoQ3x/yv+dia4NFTvelOp3VPrjkva5yl6RJ1Zm54CSaFMxmbVL6dlsoTCiQ
LAVZn/K4mywwqsjS6AD1eHR3Y73XFQiAcvfdQvlMSqHoYAqPexIz8TccydQw
9Q95LSLwpo3X8AfL3cThpGShlVFxCZERIsqa/JF9mXjmLhlibxYxOxNEzpJ2
WcdpZ8M2T1ss3ZMVuljY26DA+aFzkuLSDeJ7gTuw+rTp9bH34ha9FeRrfTx/
SfZc1xxDOwG68IhRPp9RJBRlmqQp7+L1gsJvBk+Rp/ZggNW3P2+D++ac88fW
G65kYmIl6BnqTRNxv3irOMWAHW/m77R80GwHkdooPvXHQCtBXsAuwJhAIdDH
qe4eUA0p3bVWOLGkkYqYE1vviJrVq7f5uuX/Y6zpaY17iW0p+LopFlfWqEAm
VEdRkj2Mku+mqX8V0tayM89MH6Vr148LwylkcyGGm9Q6oFE9uFA1Os6FcRml
tEtPfb+/enJXVVxVSXl9o9HKQwP9SvBrYQXsXONMPXCwmb6YI+3ePJ0P1bo8
W0q5uekMOJAKXyZjLlZFXPirFQgHVUN0ZaEZFof+x6xrhKJEi0UC+MFG2olC
phe0xBV71QrtcgCDTzNaASU/xZqbbMh104yqWdGxB3QlhyAbfhXrQiKw47ka
ntDC6Ak48uEJ2Y7C7ZzYE6MX3Lu4wfSPWAD2+ZkvwGyXDbWvtyowmAl/1s+C
3PNboZjx6qAoxP9tsMXa6fgfLJkBi+rszWOmBRLmdzY/9HtCRiaK16TjKwmx
kOQJhGO0GmEVqa68svUwuvTox73I2PgUGWNCV/+UekNdm229HnJrvdsxbnVE
CxvDXLYXPv5Lw1ugQtvu+qdFCYP5JWSyVXae4DmhBBRKZ5I+sySUKo3W11DP
anSpVOD6ctHVFFFTaeAt36dgCk+X/GrYDQfMZnYp3zb/cdhzzmwykyF5r1Uo
aWAyoCncLPRWWmT9aplxb4JxQCcDAnVXgayPT/IDynTqUPj5gePoViI5PLd8
2LFvHDlGD8IRRcxzhDM4XnBhFCImcB1F6ngEA8BneV7fo+50vD7FI71uoRCx
JBjimU7zjJ7TeXXQpyS4zANkvzao56o1V6ttHp4JGK+g28vcOBq1EJ4SysFV
Ldue5WlKOVE75kX6jhIIWb/A7L7Wyb27SdqY5BeEMqOD4U1UPXDtFiHM0Msr
rkEXIDzpR3DIA2evTPS4JK+kDYpjEVDfGnCdclGEt7tnuaj2RjbIrTsi88GG
CH+AXl1h0okxdGOBe4vh0/XxXjyl6vKHVBEwibLsvyhgrEbf0h/Z/0MTeugd
Z+KehFeH6p576fkhRoVOMd96Yk71qnHxVNgpcWIaCKCEyfnbEM16FAA+r7Z+
LSIfpFiyFQ2WiFYmV/29EkIbhKy5runFdMMyQrtTXyaqAIssDs/VHtcWp8KI
Uv1J6ntQZKMA4Hw0bIMgC0F5uLwedOAODy9QZ/TcJ+pB73T09fZ1xNCn7MhT
yeroVAkVBtdCitDOUhy0RqXMACOIAZZNK+9zM34CQPmhu6nc9IWHme5YzkYY
oXATzOfXFYXZsa90usJgH5A2hqaBujvM/ij7d2fD83K7NvEWzVTY48ohsMhc
MIONAgstXnyGs3Ehos/QXkEIegtpI7PzriuGRiwds9lnLvhJMPqXjpC/EHdZ
RXqXlTY7j+u1czi7/LMIJWwtCyDifajshPaUwcCehRecHnutSxy8yjlYWMrD
6baivVICaSrD8WmBTlJfWbMMyza+SoD3WZyOil+FqvxJVEuYlaKeMKS2Uj9G
c2eP3CjWt2/cYveSoDyt/s1g5QTHYTeGA797DgOlzkQP1hFdfUfaVgPdknm4
fFTrm1+xhcscuvRrry9V5rZLRGZAPUP0WH8NBvIoicLfhxYxRkADRyJXqcJf
iLL2Ia2VZl4BT64FWcwHYAn45XX5NR5bq8wDCFv3O/qtCmrkPfbC0Zcf2ZUf
BM6LBLnU5I7q++PCHhbSGz51ScZuELVIvtd2ptvWVRVSOyulgSMbV4e9Olku
IePD05SbRY4TssFYvdt8x7pSnDMJvoWcEUep1n9pnWbBal7uleaM+ObT47zu
eo9sCwGmeGxqi8BZag5mD3PlrGXZfXGLz/txE4aGjx7LW6BCTxWNuW31VH3M
zA2AQi0SfWVyHPpXdjz1R7iASNkX9qyyMtZeEjYOFnyrjrsf7Q6VNtmtbgIM
LmIA5OJqtwiqz7oYPGwuFWHVapsYV0otYy4jp3b/gZ+uBtLL2y08oje2DgDJ
GM8mESpbVkt9ZdVrhzYio7X3QDjn0UJxr50WT1Qqn84c2ggvfinP3lNOmR/h
wB3IAer90I5okC/H23iL/PvXEbMBNXQqIkGyWAO/qt+hxkxs23yT7vlyrBie
RBPedr2fEW9j6H+y5pxDIzxYQJyxwZHqeSRmoM9yBAf9FPurAdY3BCAZUy8a
c33RyvLxE/2O6k80gVfuVMSQJincP6wh7AY0Kn9eUUhQjao64JW9er5nzAYA
m4IdvO3LegiV9dFj3Qb4BY9VpE8RXGmOj0Uc2q3iJWYDo+1pfjx3wurWaMey
0BUtA4HJ5s4HAKOBu4QNHXaAQs+nHRESHyzV7lPl4qliXKrEytWvH2mflGy2
gqdsI84qNer0qqkg03dUUtTHA+HmXeYlDWvoZ3Tvk7M5AJcixVYkaHQesTzH
K8CHSPi/cLhqJOlzvAnsJBee4ln2AK9fZ9LGZcu2pjfgriNVyY385sg0UVJS
+R1hRSppAhGRaqeNFEZbrnx5IlBL2mjZlpfnXj/zSw+H0yMxvGzJCxIb8Bkf
luwSbX7KGYkD9MfNFk5Jo/OOPe/TlIme7ElugQh9zvUSub8qrnVxwPyYmj25
PLeroxZ+FUsa/14sQTraLhLDKvMkMrdOVJhK3xyAo8i58z22Cdyw+MrsnrTc
zmYZJnb150xM2iHLf7F3nQhkESmvGTEBt61u8INM/Is/Ei3KAfxE1L3STLr2
qe0i38DT+JKZWca2FXYK+cmNYMUrJB5MYXw4xQX2iE5mRTNld3dw891jSLH2
P4O6NTZ3Y1WyuMw7ICcwnoAffsqXVr2olsj+SxE41UbjzceR0arnGvnNSrV4
P9r6SenV+C5r/vV+djARRNpovKxynZ/zDgfkd94ZNLkM4abLaAfJlISf45No
Di0lqAhhZbOZ1p8Os0YDKSeLmW782PURd9dVgbzXW2e89F0/Fi9E2TzBnke3
JuI7vnbAN125wFAlLRJf01J9TCsEs2zq7/CLtZNiAaRHLYXiw3lIChoUVMv+
RF644CReX30W3sbpC3J/0T5q6c5VF+Q+HCQYH83LAVdUimTqIGf18DH6DGaM
l7dd1DFpVLZW6nG1Dgu31fZQsNJxCd4iqFb78OJK3r7DKfPm48LAEL+2K76r
IzDCNEI5KKJmnn+qxYYpayjkT6fI9IsEk6kwze5+lY0jGN1JmgD1PRJo7DE9
bQEsrFQLAmnW3xLaI+DrpMkF5GxOsK2auIZHoshdEe85SnohcIaqzn6qyFBg
278uqPqhkMoBQljxVsdn68f7ZEKsaDbkFdH2fGXn1o+EqaU/zgCjKzs3jclz
CClWyZQmuVN2Bu1jVt3E8dldN9QC7GsF+ESnoICijuX1S/V2LzyAEt5NARD9
vz7CfupNlLUpkmZjYqbJKXwwyjAQ5CQ9WK6hqk6AMij4SxhWbgHFzyGJrpZJ
3zVaePoKzmdMR1G16weBOe+CfrpnGRcX7VdQlHF+LY/p71DWzDAtfezOBhbW
vwV6qskOoXq8jrS5DByrMD6KJ2Nm7299QiHMFfd+vno7Yg6z2M2d1T6VtLHT
qYeA5DJ1PWRQv1CLFgZo81C9oUB1C9glbrdz++pUswa7rUdofaH6Te0s4K2B
ZuFBP/YWivnplRo+GKnVYWdksEtI/jUc/JnhZsJaICwlpIZ94L+S05VlzaNF
fZTVAj3VIEdIx22FkWj2umi5CN5xGccPpl0x33uekfGn43hJd01cxZlxon33
rM7ppc0OX9grR0FSOzaTi6UOUQYJ8RoAD4V8A7aLN4YrNMD/IdbNezUvKL2t
LeT+XJCezcE7Wuf/0rk8xD/HdxK2vsLnGkk7AZNsHelNsi1l45PFs8DL13c8
XO2T1K/VJA/vzoNJQdMw5PvuGCSzwqQ6en1aNkFJ/0Sx/j9QvaiGGmx0SGHM
eGuYfNAhMUZw0zA6yDnQnjTel8oeO23Ffzqgk2v1/Vd+/El9v87egwvbazHu
7ryx6o6l5zTBLuwenH5IIiPBpHOs9EauRgY7/BqMbRWsj37tYPKzH1mzKAiU
XOcvkplwpX85vAg8aBGUSazGaPV2tXNxfzox+67WH8Sua8OzK4i/VEFNE720
MuKTq8Oax+VMc+GyCi9/KCaRXp6BA6M+Emuv6fXSNA9rnyjsd1kYvPCpmUY2
ookb9kXzambsq7Bw5bMx0kmRTeKni9LjwzXKBSyDzcKlOgKrIvgNYVaneQk5
KUXzOc6LDZNZOMuX1jPrqkxSYV/q7PeRH8XKqrzY4FR9jM+5PEd/T2bhzjb7
q/4M5aSM5gY9v1XXG6fuaad/gcqW0iFgzyjyJ0mJeMelit0eE2tiJAi5c2vt
lrXbdY1uEKy1QEGR1Rra1fHji94j5s5CXvbmRZMEiK5sADKsnMw3Fr/7uyim
SQLV+RU5KRHYJEelddmeDybtWh6Pi79p3V2y0yGlZfdgMrb8HDayrLrui0qs
dUF/N3S+rdxyvmp6uuzhtBMJokrGj14wO1R6CAuM0KV9yIxi6vdBiDOTMfMo
g8NT5+83GJZA5YahYaBwNnSv+3V5tIXAEr1dBEm3XgsI8N8G81U2nML51YOw
ol12fs4yjfIuGcwReYrfspk1xt7BnGjISvHcqHKJ7n+YxQ8jQYYkMSEa937Z
x/n6fF0amk2tKTnYeVoTuR2yAgFkqHmk4icfb3UqFO4Xf5x78q8FIuLZUhAl
JK2AMS6gGNIWqz83rlKkJZpc7QZElZfTuzF86Mi2wYuQ0aMIr11TsQMfIjl1
Q1b/G6mspk8S4vvqxLI04WBlK6sXFpNbbj2a19Lew5+XjQELDQvKzcCf9FCw
YOdjEzuSzbFSj6E3VIaD6hJtfDc16zkW37BWDDuTo/ZBhlxZwXm3aiBlaoMf
Oz+P6XEFQF+Uppdadtto3FPSovjPfaJZAjnySJ3G/+QwKbg0anX4bAGgmHp0
PG4Lgo4LS/4pB6hcdw2Y4rrAL4EUvI8dn5gpJU/z+lhvz8Ux5XytrlXXB6ax
bkNuFp0IA03QLEkLjg1ff5wH3P4II3mozfVgHjrD15aSPZLpx+kUWGJKs+Lu
BFL6ZLsVWCWCo+B47fZE1LKshZmxybzRSAjlMw6BcO5mvHWqzy/znm33Yrdw
qhzxcb9R2LVcoSyYPO2KvDRTurz775fZ77QqtDw+bAWoaiHym7+2cbC9aIop
SAZw2YUjo8P8hV65NSE8P6GVo4B8h99+NTuJoRknWPfD8UZzJ4Njanqk/djs
sAn+gLUzzjBuS0/0RxGrHsYa1crZpr+0w6deyqbjjlNcHa2LDmrEl7REHY/H
r56x2cw+U0jghlheW9p/eclAOiUGX4ygZxEm80jf2U558cZKhS72UK1SwAEF
/YF6YNKLX6CYkNUDbmlRVjEq2gr2671e6OP9DWKJCfS25pZPusuuZL9M9H6i
xgKfKLyUVt8P3L0dPDjNAAopZwnEqqvehyb+aV7Ifu5wZWEk+vHUdMiNcWCj
T2GShTNh4M1c1ZuxU6d89SMaDlUO0PIl0Z+STC09h/YLOvxSWY2/iaTWRLrQ
PCI6ZhnR9370Pr2o9o/TwjvlYKI7SE3jaCyk8HldisfZk2RR4z4qTcljdHyc
8Ujg7Hv8raDQIx9tR7JQTBFAUAHvpY4kLzxmuYNU8oc30XF0l4YbdOD+Hk91
47/TACfim5mqcQH1b1DOsQs6hm6ZP0y6PWZkuUsfA33M8CGYYQdvQsXQgK7c
TUszC89rtjey7o0qb8gPamWIzHCS05WX2TljRB0S/uoekejdJwoUs6weX343
1/MuttlNytvrs5moxdgDdiXlyF7aBQ3a9BRT+OeOt4DIupjr6Wc1giBZOqVK
9LhusslN4TKANQsdiWnAI9RKbOVKWQX49S3v72/VyvMZA/lhOoN6X3LVB81T
BXvlwYhjHLuqcdqhfHCzVLNTrh9CEBEpAcsXUskwwPkxwvcaMmoBzxGPyWQH
BZCjhrc/zoWRGBsXn+ImXyuz5b3hHVZttTqqrHH7PTD/e1iku9TDX5X72CK0
2JPe+/8qjg2qzRPZuG1Mgxz+QLGUDxHfppjZY42Jg0TJ/IXcjOEzjitSBBYN
N8rV53ZtXtlW5qX6TDaNMKCRdvEmT/a3M7BMaXIE651ROZqk2xuPfObvIFXd
OFy99hTvtL1cTF05lphk4I0+AS36Loysvj4KH4IZrQPYOIh+DCZVDtuSxpO7
EAg9HFHa8hnL5WCGOM5RbKrR/vXmk9RHqoTKpo8cn+TrZrWfnBl+dXRyPXPS
RWlWQYgFSfEVWpXswRcVJMd9uHngUjhP9nPv1Dl0WEfFsuGQfpoFpYh2UtL/
9duZ1wW8WammuChUVsTsAWngNdyNQMWBABS8hmhl7eH5pKibYf6citR/T8wf
gL9+rZHyVp4pputW+q0ZBFhZKbAB5Unnw45j2cSKCkhVwRodlgvuTZYtsaVH
yoO8kJIgw/bDLuy/02hcGBBu/MwNl1t2sJpB3AMIPWMTuPXcKNkm0jfXePxe
RsaX/TflQME2HPwK0rOak2C2b8AhARPix8UcuJDOaLd4SrV4B9M0Hx/4UFpt
mj43Yy4Y+oigrXxQOmC8CafJ/2Ibpow+hXprX3qHAKWoX3JVqWHlz7gtGo2L
dR39BOx7USaOmzmw2jKhx6e/uPBv/2Day5U8iKK6O2nNtmgrsN7q2+S8w4Db
wlQMVS0O/x5F0FtN8U2h1IqYGUU2COPqt9loZ672d19eL4+jtIIOa/x3uUm6
ejMNgy5cP9QVHa01ZGrFGzVUKbZqn5SGtHOt127EMNd2XuIObJ0pHjX3Jo48
N2TQRVyf9/PMepR5R6vH/GX9KiN896tECs3ShpP2J6kC3NuhRUKJ1KAxa4Zk
drJvEhSxMeTEfEfDy7f+WC/1KILg1uAvB0M91mP17gYIhV42Y3HEHBtGHVb4
MnYJLvD/sU2CCJ+gBCdZAqme8BF/ryW8RJpz7+6ma+c3lctYvsXa5JFBBX3D
e2j0JefN/aMuUFXXlEwzpbtK6u4UqboA+DMG92+FnxpWYRiwdQZLwcSTfiYv
WWXxMpfq3Qhs65dAZh3Q3Z3yrWuIqp422X8Y+LIxySdWHmHZFcaMFwYY9qZ2
WNmUFXv3CLQODKYerycbBb1roHkUAeM2nCeCrKHI7SokDbLmKOGaSYm4L+QE
K1MJe/BLFjTWD2VaV4MNOvRCztHt84PxVupGkBP3iOJvPiysOc/VL2DN2nJt
7iGOtp9EiHNBdr2KuxCtOxfIEpwgpLl+xaCc40AzpAjEVwDWT4y8FdRIUBvM
eG8ML9lNl2h2Mi8Lt1wZ8BCSLaSGCUmS6m4XlP6w7GwfjIZHB3eLr7S72n3k
ZSaTGLc66L2SJNFMmbWhu2s/b9wPdkGcgL+ydqwdoz/m/8NN6i81c2FAHdrj
heyOwzWtidmVaGoN06XUdSo8GGM/Tjc2YCknCq5++gmynbG9D9vv+fY5iGTQ
XoPNWJkz2xEWbvqAkkLuqC6p0Au7xRPDaXSZ/+mT6wnQ60o6u7zPu7ghDTh2
jJqrNo7LJX51elFHy1/Rc9QZz2YDWzQYXUIvsaDVl/9+p0BJbLRGfby6yK5Y
/UYesrKRVbB+hC8wm/7asgckwR1oT1dsn/ImkB2+XzcGKYDYBSIAN/vZyBV/
mnRd4YItgybXUFfnb6K7RabDmPouaYEd9xpE2rS28xTIGG15yzRuUrqCWp9S
yCkWFdKPSD+tLjCmZMadR2T1VIssuQfeZmg1ZJtgjPwpjBInhpb1AW+kn/zy
JW77ktYo2udWiBkzlniUjoqifCSFt5VWKSxOhQGtLb8f8nWeb0G7WKcozIWs
3qgtjSgLm6mgNt0QgXsBofnCl8yNMZstXo7hrEurvQf/G1/V6c5CHcb4UbNi
7HdjZgUKncpCw8Lil9eKtzq36XU5uXU52KVsc19re1x/8JJlwWngIw5OK04K
2mjGsEOAIznj6TLmqdtZkNLRbDD2OYUlbg7jH+g+pBrV77hLebFtj7rfhWZJ
o9+/EP6QQECAjYZWv6bOAcqNhFJx+bs3geq+f+6Cak0Mw7pjEbWN8Y4huoso
BhMYBlXd1zsMJC1Xdzoz8+HJsWbjzTpYp1G1+Tl6AaSci9ov/PhxdBkag77C
6gGcGqUFCgGit/0uqfi1VfXhcQV94VZ0+Moj8aHr6zJdg3yzDt4/HacFEMh9
D92tcOh5CBavuffGeVRLPtZaDGuYXD4+TWlemTsOr6LGH8/Z89VuCbFPde1s
I1NHTEJL61/JVyb+tcX6ewqV8CgvZbHqFUSvfgwBNcq9R8JsPMGnW6/seZJd
E5vwK6Df4diAUYB0pSOvxBwCdNSCsMWhcJA8Ei75SIRgz77OJrQcm8RGdwi9
rnCA1pqNaKpXc3Q+QrZ2KNS6WBrH7d8rSUssDg9eTsU0R7RB8DnUwl+x/SQ2
lTOpW0ChdtuP4HywY+0XfWxy+1vDGwE4YbAKXEoNGY9hTbqs7bHdgWrVbXNS
nJZsfnM03wU+KyEKJ9g/BPzE0CJmt1/bUfpNnGIXMIheVI9a9QKjURndvBTY
7FugahEhhQ4feP/gisuxsBGSbVrzShP6TQlYYOybRaMpwn1TsZeCh3QwreMj
PcyCuxLbHohnt8E17Kh+J96uoqPUmrdQsv2CIu/ntdjC5TpS8Cks3PuPAzkT
vkvY3aN2PLFezAxFvtxkfL8J+fDg2WEZsd2xp912kNjwPs2QqZuFC20LaXdn
faBv3pucLFz8/OA0Ch0r9VgP6OAwGmT4ej1fiBdEEiJzDCO3wYvo5pch3mvl
mTH4q73u3DpYzrwGtTxu3FT1R+A+e6MDhrb8qPhFU/tMbvWDEz+ycCH2FfrD
QrklZKzc30eYJQkXtud9mTUrpWtR5WAZ8KxjTDLS1oYWqsxqmN+4u3wC71i1
TC9mJ3F2QmV4vZONIc2L0qHkxXibEi0EaBmbLUgh0RONQtse8kYcfTTElxjA
8XcicXs/+8lMkZHvHnRbaOEYkRaY0yOhDgC55VpH7V1AYXXnxwogH4p0iPr4
NFWLfPsmKsBXn5UuO4aW41ExsUDs4r4hsZSV7CTP8GKMl1lr0woofvJIpOrF
Dq+zcTzE5tJ51SHkhe/pb3j+a6pZE5QWtrPTlFFLBRHbws2ZSzeISgWfxgs8
rUQ7dYmGDW45fI5Kox8jhE1/V3f1g755J24a7DnSdY30pJeq51c+neryVz7n
5evyHOf09NGG5OLbEhC4QPfP5G0qcK3vCg61I80X3tFdpvB/HXQD2s3vD+o0
0QYBk00Svm0lMWFAB7nVbDaBE+DTRp8Aj0bIZa/TWsv3Mgms2oQICsYQt9ZC
4BUMfT34OSSo4rWMyhldIbJXoNIUpSeihgnZLxnuZC3pZ60rx3PwbLHFdoyk
Xb6Ej/pbfKkMdhZnpnFgK/2kbxEEFXR3Qem/svr63xmr1jiMwp83JYJwTmnf
AEG6AcPf37suzu+XYKHbnKlidU5Rzq4oC7W8Sr0XuP2PaV71zpwawlFr58Xr
y6/Cw+CNRURSqP2mqL+IZQHt2kEBeb4QWR98SYu6bC6aMLA+tdnRQqbqjCRM
pOJ+edpwEIQwazXnSL3spTrDA94xh1LXrssxRdwEC2QsfephRu+VuV6/pWrF
MSR6KAxzIi8KycvWrAcJsylDEUNIQ0Lz74Y15ptkz1WkG/M19pESlTqswW6A
ritZW+xQ2NQ49HHNREAjU0r9V4T8AbTdqb2lrCb5xOKIOiyzqmbS4+6IDBCq
HLwjDdb0+NQsR3e8mLoZwZeR8zX6zG8HUlY9SkI0/5M54CD1eduuCOVy7oC+
XZJt4F7M/4XW+hT7Zpt8ZMi60g1gMrB+4xb13xRUBUP7tzBLRL6UBkWWENss
mAFu6TRhlnhNkrDeL5GrMQOPHnD6W8mS+YdOoE6Rfld+/tqxr8fJO8PB5WdS
uOK8ydi6pTxfNxcrk8ps6vpBFIHfDhfFJ3LJVrsoV5kEqB+HKbwgM0caktGN
p06NEVjnRa14rof2BSOsgo5v2V100ZgXig7Pe52pr2cuiMWMbZskDVDDUQYX
Diz+b79mDhpRnk2NBXDnr2JP2gV+SfJTIBjfk8uanBzLTpkLdwyf35WkWKM8
6KnA2D/RrtByEYg1T3DYnVo+saigGd5eV1ClNdxxHLWPMLhwUjlrg/V9KByu
LzCpdl72Z6qFrS0+dhrQr2RCR0kFv/kRIgzsOqQeBv+ab1kwPqBuhxDh0hS7
dIhgwYw+RwE8edDBqaLgaxykTkhDP/WXsx31To3wZEFeFXqzN/mnluohqwsy
Fzy0063thAhZ9bxlNNakWw3giglfPQca1ZDx+SxbFqYnk+NCeH9IRxeQgWkz
WUhdjEAXoUxAGUXl6b1a/OEe3EmFpZS6RaYcxSEIxd2ANiDBu/K0JRW2iMbr
djsQijMIIGPfg4ZNimHnKYByZZHkp3RXAqwVrfigkuwWC53RF3beUtadcRPt
6V7iezBHpTYbzjmej/KsjIhC733pzgF0xENGRe9WGEBea45OdEHZBLaJBBGX
2gPVlmBiaJqB/kbBXkw0cSESyrH3qSJdL9zc3X5D/M4l6c6pm7o0KZOonWWa
VegeA7zMeqv6Zd8QFVTDEQiVsr3coXftxgLW+yPixwMRkizJP0xa/PcbLa6v
ciIOCPk5S9tipAE39LJLteG2K/QRAqUaqWttZQkLtyMKOdX5iKYQBm7QqCL6
Uof6fqEkKXVbb1dfOJScsdh37un7VSVQ0akmc9HruH1tVu6vphaEHSE8KAE2
CHFuMCBCbnjnMyeqvjYWZ4+lODcjkqlRQRLEsF5XiwKolebBulu2pLR5s1tw
6jGWluqmV9smESSY6hWyHbbLV1wWbhsWlKhJjSCQvEZuPBImrupudK1ffaSE
wbWYgZqb7Ekx3TbmChDjgJWbXZjRwf1SuSZ3EXfc1zWPCF0owj9byvQqYJxt
kIFASwM4HFWsjxBM+3y58+DkU7zvjTL4DQV/KlveiFXM9kKoW4l+jzSPWiUF
Tgd5V17klDc4vXpnpRJVqJ4G+d/zOeTsJ37m56PKHbf2+P9vAetfMKLPZfF8
FbVGYl3VMbtJoh8E5jpKpuDuAjTN8lKJwNV4vUdy9G25lFcCsSJRZ10YnPKs
5Olfd4hzsd/lWw3jkUsJWE16B9CnSNwJSzhCE+yWu0PMk+ViRJzWbXPn0tmj
KWkn71si+u0cD7wf57HYuOBGjjxM22KlMhNw/XqlfFZ3wb+O4CmQazRLZFgt
tCiNvYbNGAsZNJxMRM0BEy+NUwthKUJhegyztzrEks9PakuIZMZcvyOxP49V
q/hS8FF0aPvB8hTLPWD/OQ3Bb9qv8FGckQ/DujEs50GeoCzhBMieQSQ9YC6S
3ab9WrgWydcW9o6VOUojKSM/MZG8ad+bgrPc9SP27/687LZ+YTqPdhho9N4q
+g0+5nRQSiy2blfvRpBV/HnwNnA2xzbawY0jLwQ9+a1gMpA8q3sL9+JOVoOw
iEoCjrMtBHmh+8xYX90gswaRpHII3iI4KdZj00XY3MLBEH/EoqYvFREDLn2i
3KDZ2hY/kuK3nBM5/Apu4UPhuUD3AvUYfVxm2dRwqJ73hQ/E8VPsLFj2Lf19
otMe15eiK/EJZSPchHCwomGKkRUJUJflhis56QdHFCiFV3bOceT3AJqtDrHC
8j52LV6HPIzsTPUlWxZx7FWJNzc6bJUrUzd+elIhZtcQdLYB3oIOaTVc3BPK
cP4XwM0QLE478jtyA+pbSYfxULq1hRvtmNmbNChvd9chn+P4cx6WAupAR/2H
899sFtkJf8Hff9vYOK0hggy8hRv6m6xl4pEXM2tvgXoz9OEIZTXPWdl/6i9O
ErUwKaHInFFtMaHjromeE7Nv74Mh+RhnH//8dggkQzDEXrR4dKa0+A/qL9UW
p36auwk1xF8QSOvXjrF9jQhAkgF4yuadXlQH0V50webS1hooPGOvtoZm/8su
6nNyDAsr7FAvS7lKW38ZQoHCbICJ6IcQ6tOQuopqgZpF5WBVChjKSYkPRBnB
MkyqaRfPpuYgM/8edbgemU0ZLl4pbOfjh6xVcMVCuc4Rz2ISkh39SYn4xoRa
B6q2CoKSBd5g5Jdwgn9BSjkMpn65ohgBPlcSeULiMLRpJXAvcNF5abN3AWlK
7uDIy7SKNuYYz+FBSUqKPr1wOoDQ7OwR2J9j7wVFyCmoXUC5+gagnaeXbI2l
jDoNNpo0FXpaQGeFsaaSoLxqUmbW14HwY4muoIUuLjSXXOHcv8povEDexKT8
53JzdQhCrLauAGeb2vScn6KAFpxWUyOlRC1xHUwPlb0rHNYbvxO67iyEWMh+
0yzv/KYsPYGOCDnEVATM6EcW0kyUvIvTMJw6gj2688ERc3b47bSqGXHUmnd+
+AqfaTW2nWOO3PpuZNTmOlv32IS7iWU5Bx99L8K0JS5LBEIiYF9c/xfJ075G
09R6470un9cDPXLcXCUvkGcCIUz1iGElNkNXqsCP/biGpo8GiOPdT6rlXznC
KBdVwkNk/AwA2KxOwXJZ1wP/1ze0HwdRd6gUifDvS1asNq+pakcBKC1a7h55
CDBpQQWkj4yLCPWiluwTrp+8p4vSTiVg3XJcz93OpZxg0MEv8l54QzfUV8pI
5uvuWIQW3UqPHHOkoviNQRdn1Zx9xc4WXm6/A7tNlLdx6wPAuPgYkhK3kdCC
jy8K0SKB6ZfHoJqr5NMSqKrD/7Q5jOG/S+eQQuu2SqQ0bK9lsih2ZgA5K6Du
fv642FonWpC9S2IjxU4G40xBe8BtDNbw7enS937v7GNfX7u1OpY+WWUCOS6K
TD1AeyYgyDaG/Uqw2xNsM1Toa34ryUjJO/Iphmf0QcJSLf/SyzG1VQw2IRWG
LZLm/CZX9zCwqPN2XrenT8hWmrf/kVQBtK/v0XWx/u5Pch9+PAKQLTPxn/L4
jbM+vM7YQJHsBWgJ5dndspnV36fXgQ/XcE68IUQDdffiqx4j7gAh+CgSFE6C
KYklC1kxDmDymRjw4Erj1rn3ftPfJ7M9V50eIKNbrdCHDOZHXXmNPsv9Ur2/
+hM9Ae5TLZmg0S40Lz6TSPscqS0STqcQdpXHdeR0u3THZX/+RGSflBOAOROB
CCuptQwgDi7iwbn4a4wfl2ju/KhqwFfrgOlGu3y0o6DdYfji71j7mrkxe7XV
Tb/I+pSUoXWm+dvpbh99XjCSX8JBfiPwHCO3kFqfVZ9Sd7mf2eg8iYKf3ZLs
dzb95BpL913/N9w5XOrUtyyPMcRMbJl2IE/eUTBhoML6TNW0h9XlnvSLkHNa
PnwqZKY7fZz9Ioc1qmO4eMAZxX1meuzzZqTR+QHmXzhJEGVPhfDBZIGOs0Gs
tttcJ1uYDd5VLRByjOqDGEeRXAOK5Msq/TyVIqKN8L/Bq44Lu4b0SBQfXqvg
WHLa4jwVArr87ubM18hoI55G10oa3b78dNyLgmgkVyMzqUGULTkrElZHyPgw
Mhf44SSNHrlL+ZVPD+z1efee4Ms+flgyt8aOVrMo7e0SHrwapyaIqTfxsyxB
rQCfDrS9OVSQhITtv9U13XFUcTTJXTG9gAJI5yRYWnxtKq+Puo9PDyGc1O/R
TXq2K2D01CdW9GzeMW8D7wMZpwj7N//3BwixVZ9d3vWFvh2DjN4cZspbmmB4
FWOwLbmMFvnJB7d5T1YeK6v7ODxknZxiwX5SXTzg/AI3INMdc1t1Voi6UJjT
n59TADzJoNPRuvjxQvN6P3IoPK76n8W/G+HcBPJ3e6OsBYMRGRWvzQBC4hf7
F1qyjaEm7l3FDEnl4jnNxAojWYQBhS2vuQLeN3zK/IjJAnc5A7Vmk5AOidUj
POcu0PzzD/wKe5C/wTLYMi/1yuoPCSmGOT9M97qQ6i+DCvK37Mj4JcCt0JCq
vU7sDYMLOWRBn9MmCtF5dnpKhyp9FZTg7JcmjApXQs3CZSeq1UXzehZb6kv8
btXWnvWFxHL8JuyjpMMgChc9LJ7Yb7TUVAHgEx72jnEgni18jSCNfblpn0oU
fJ084sjdHGD15oLGSaSMAlCcN3+9G7dwS2p+yH3l0xgPzc47dNG1actqLoac
CM9gDU2AK/LHHLL175Gbh/QVtypkrrWTnW6zEEG1mt5atgctMJBFVvL7fJx4
yMEQyaSeHCd+0hHo5qn+grMQcXSgyxpBXiyzRVtvls+Cp/yXoskP2O0aF0s6
xyZ1pAqcIDIxO854WNE9XkM82e3tkhOz5Osxylm5VtPkfcuMc3hvjC9kXMI1
5k/po2VZRAlYUg5NGpFPPqpLQMk6EsKsq0tsJzoWpTXa/WsRJqLnzWtrZ17m
GhopkWQW7hwMXu0MDNzxbXrRawf+76GvdHa8bPbTQD/yckse/qDH7ohetgBw
J7U=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2PBBpLod9UKG06DRjX3P/TSwXIjVo9+twQ1DJA6mrlJp7YG5gvEl3ebODARMkFBp7CtxNrtgtMi8KyP03UwV4hwXPS6ueO9H4o9OHAbf/S1Q9PtGujpeJJdy761LDlB6BlgWC+sP6skesRra8AeTmm6PGsOaG6ay/cukGRrcFjxq8LdKdOPnd3vmXnPGcr9utbXQxGKw4dfPtGcQM8pr8KiVyQev/ObkrhJg1czolZp8oig+vI0xConKwdxwzxfr6F1UhstGWOIUJFUV1Aox/qfv6sePt6zwL/Yk+/vZlXrjFOXrsMyzS8jRtxgTqg0K9XE47ljPpvigk/DVT7t7Z2ENCrFJOiUNEf7EKDn0Qevpo5V8lRToKTjnjHitTD78/j9bPmbydw9tQysBaZ4a7xBOFm8/PAGYetLr8B1EwbN8vdbFecXjXvkjJV7apgbzN+8y5sNJ0NgrhYqczgSz9Zpn8S4ScnQ6DtIcyHAhsZoqvED3jVakjaFGm1fexKsWFu/SMO4G4HUJMX5mcXm3QHGLZpPh0i0MiQxib8ihzvcCJSAgKQhFibD25pzsebUHMMMLf8NKVdrUpAMnoE+rOHunqkmSTd79rwqUuWs3s8SFP7Su8rAvfFwCHwwnGY35Xj7PzM8iHxPhIHu3bswI//SgRub/2QZlZyGJ22YdubdoIYa32Qp5FFz9kPX1hRr4wQdYwmXB59sxPzkT6Ukfo8VM8dggOy+kj1jFBP5Lq5n69mSjsodwXDTtHhka64EgDejGTF9jv4GMLcIFVag25tScCC070FIL9sO7fxfsuYxdNBHpopZsiEXZqwMbkEmfdMbaFoNG2QSN7+cYiPlckIspIMCVxHaLb6vgonlzq8mVhAwWBSk2zPbIPdgjJJnbzgZWnmZBw4bSPrppCjtK9Dat6gjI4QzNIu1p8UYGwBxK6zguZZgzXcrbiy2B+aZ1t0JzjXnDPd7UhYqK6KY09T0EDPBHWZHXN/YJXyAuPyyzJslc+wLDCX6RpZXIj41F"
`endif

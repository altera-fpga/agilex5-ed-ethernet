//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ldQ/JjNxHgz+KdeFcpJVD4SffwpQi7lCqCp8Ynpqj7CHLyLwZwrdZA+wyr8o
obZBxwmehmmIZOh3x5+TuPWnIX02X8qfMRnPff7tnQJC2vOuehCqJZDZbJBV
xYz2+UtcFBCfRwnCzNyIKcBsgl5SIaCxSxdwj9xr3uImE1U1XM+uo/jvVRbQ
WFeFc1jnLjX8wRDElVdue8PehEJLZ5ghqaqxARIVKmQVrAf9Fid2Bf+4lyPs
FB0HcIKrwP9BehJdxeq13z7ZbHDszHQRvriMD3tnSi/zgiwuNbx+BqLC490Y
opeuu0Bm+CJZ0ul/8iAdJT4K4o5gsLrtcgWAyaVFJQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RXiF6muY63UHjwnlwBbjOv9O2qSMs5Us2DSoJkm70c4I65lD77hp0OY3JfP2
J/b0t8ABOZV+3TGzb1pZzoMF7iF6wHXEkRDQCUtDn3479wetpzoYycejXFlo
JFT8QwpLlUSVi03aZHibZnZkXXK9wrsSNfrmCAsXJLIOQq/URwvAgJUDyA3d
WZaqSjgl5d6vhISxXa54fanpqJzauBgc+lOkVRx80pmSgsCymYHCmmbPH49E
5awaV6cavvJiGI84IOuAwOObYnLJlIDcMdJ9QqqVwIuvXVxOQSe3ZzlWY08q
fRsZtpW7W2goXqEmRrOLtDX3Rvb/0p6wd0eRUBoK2Q==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lM1I5/HbeH+pamEtVh7y5qQ0xNKOWqYF1diov8Td6Wgwid9iB+iyi+HnD873
pUIFdFVQqt++aH/ZUCMPkS+tVIFHEKmeK/BextpWPVaCjqtLY5gVzZYzbJps
bFGMv5WRchyvoUCJ9bmtfBySJg8D5qW3WW/OmrWLfo/4ed49TtyzFDQy/HIZ
zyrdn24gf7HDZ2vv5pdEDhmwkzFsse+Ds3P1xVoTkPOkpTezuH7xjXkJ/lyn
1mrFMbMu0gGcJ0ZPPTZbAz68M6rg7fAif6hDG/O8Ei+b4m2UZbhCuo/Dy+9n
AT3AC8BLhqS4A5iSQrUZTrUrVLLSpWt+ypPY4npaCw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G8CLdZNnm6y1HHNyiu/YDj0RPnCXb+W6diCsRiGNj80KoCfctLpyRmjcMBdW
IkDXfFVN0pwAQoR6X44Ont6K6rl2MOg+WtYrP1kABKJvoZwL87c3tnD99AHM
T2JjCZz8mtsWO93nvFmeQg88YRCDB3svUTnbQV81A2Yw9O/Ax+zV+rG759wQ
OZZ2/C3dsQadQBRFMrJpB+U52Aox2gOacNdWkYPtHlgHFgsCIE1aSDb6HBJx
xJ+w9obh4nAxVO0cGxC6XPSMLVWYTMvkItgs9q1ux6jyPPVLlvDBcxPwMMRf
nfW+Z9ge0YOpty//1H5GYJlH7PdvSLn8ynHNfMU97Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WX5YI82fetc475tOYb5G57PPAklia5/4GW9+sIQdnJ5BgstTTPVTrvy1n1VP
SP1eledjgFFU/3V7+5dMRLPVZ6GyG8dL82X4crnN4uFxSNgQq2o5SACq693z
mPJ7ghQEhM+3WM8odCJUd0hUWSCWbi3zg2dqrM248SUI1kMbTqc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
likXWqA6VmsrxLcX5GbDTi3JO48xR2bXhGN8bHy/pwgdruLlO3NoJzXBcqRL
wPYb/nLFYzkecbG0iHoIWPFPmRytZ2oGDaZOs+YR1/e1BT5PQs7nNOjbPWMP
ZemGnWPwDmgd26d56aAC1h0Q2xJzssXA63Tcubj0LX+kR31V/DV4EI/iYwI0
cVl86y2acpbzDKddXoM8EskLg0seifXBqZcmpfofV4LRAfkXrFxR7n8i1ke5
UEBvGKExXKHL6zwt/U1VWMaoAMjy+0ok1e7mjOep/xcgHjZO7t7CL3dZl1VR
ox6zP25/V2mT7G8RCPh5L3n/J5I8+6wDlmBzqip5vNn3swqdbSCNTNUxpdnG
xyDm4+tyFdrBylyl2HEnCIYD2QDkkHaI3K7GZ4flLavjOnrjazJ0DfkQjODB
wWHl9fnURcfYav7jtSpTs2zj+0YUcCI2LP1Lr2BGqX7BAZE1ZGVV95fAdl+A
2UJylRknd2o0aS9kwACG1rHo0sj5oubP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dRpRmbw8c2ypqU82QiVEmwwCYM6ka6ksK+qP4bdy47VHL47XwwV/Tj0Skk+e
CuJy7QHDM2OKAPaquSjdMscR6scxjh+gxZi0UhCuj/wVznc7KRtjIuOag1VA
mqVjqIfWyvIqKcCzzlUZu3pf+vuTFbfdkbQopsgCqAcAfk479eo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H4kZuQVLahv+iWi/SlK9BHkI7AyC+wNcrPS9ykySXn2voTdh1efGd4CGBUgF
2MIep4/Qn4l4NZq9lEbLein/9ZF9hAPBnSMMX9Ebk5PXSLCACJPZIJijd3jC
SDq7vKusg8lbS3DamfSwgiggaAbNkrH8a96GxeEeTybkJzLlKLM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3888)
`pragma protect data_block
k4IZNFnKZJAH+ft9XvWide3NdoynPWzFTtdFIZGFhrHT/AO3j6MFnOhQ3CPM
PBub84NnQbAAXEebkE6OjTTrVmw0E18pWXLH/Wry3TPz51Xju1HJc1lniVU2
oRDTHaheP9Kf5s63i1hjSq7r/SkD00ZXeWUqs+Tm06VGUaauXV5ntE7Yhz8t
/9YT+KFWIILxrF9C6fc1S5PN+FZQav/Avwh02mvVv9dnnx7rpZgTuZfbfmpl
jikiVA6jycvUTc6axvOjq8Ed7ojH/JyVI9EOSn/SIKST8xP0RwdIoedSFRQ7
RNYtspx1vBb/gkfO1FPNv70JM1AWXOHbth4ARl4bw9DVVKnujVQ3pfP6v5gA
rxkd5+cXFVHRJjuFGPFdghTSdrWKarsOGlEAL39tZJKLZuIjxlnUEZiIJppg
R3njf84PTPMQCoEBg6lyCue05jiEIJLtT4RPF/yn9U/rUkZZtv5mIsCb/YAa
Yv/Nx/WGJGcwh9EK9BDfqWxMhyQbFB+TruJHKKj4nuP171ZG5B+ykhKaCihM
ZgAEc7KtunSPsvBuYmCMbeMoH1Wp3Z4p46oBd0zUIE9qY55hw/a01tkMDCIq
yAF5zwykfoQ6Da/h894jFcitneMjrVJZL0Y1uI4nZd1Tx0HLcMZ6oKvsT6Ju
pgEghYIRZZEAfqddaLxDvQtnM0CZQxQOosdP9QY8fd0E6IefRqmBjTSrLdoC
jIL3MuSZ8lixd5eVotZ0Z1JiAIpIb+N66t17NYC85Ai005Gy3Qs+n87vDOqT
tyIErbDT6OJLa57hN2IBeJ+ySHKkkbxT9H1k1+xw2RhXF+t/Z1wE3vCgNv32
zqu4BP0iD56i5VRwApjJ3ACOSZoqY0TtB3Te1Xx8c736r2o+WIsygf8d7iVC
UfMM3hPEc5jhvUsIixmwy/7WliToEuTombfW/nyWWKlu11J2UYvuWwK4p6sr
+SzIYK9SgRyoZJM1GPsS5Ke2ulngBpXdDVaxx3UwYlzzsu/muh+zwK62yuWI
Smm9h0D2lgQrGk2nB7LMAOrVPyiGzkAYO8n4VEllvixZ1DVPmQpCO/jSRj06
MtFczeyMR/9R6p4qbegCjR1mnV1b9XdIc7hEA+3oWFPpJw+sCedNNeaVgvWX
vhmg3Ivv4gDOZsixMM4mTXw/exl4Ynhsu6DTK0gngszMpxysQJs32J+hAxDZ
0LVqQaK9vV67qpo84/57OC57UcnPkvizHhSoqU+ZCxGX8uVIadtTrJUm8o4w
QVE6m3rvRIwCWqwjALzfMAFaWJGp+wOGniFlWszZr7vyvVKlj4CKdIbWiZyU
inJ69b0I+ybxd1OzKCPLYVIwai0PpEu395h0cOGUMvT2P1PDfnXS9t3uh9hD
J7FNyX0hkC25G3E6KWQ7ze1REcTqz97ocTxIwB5ch5VyFlexSE+hhi4frtf4
zFQZAgozu5WqiONda2dxrhRJKMosg1ylVeGtFHiibGBmNyfBb2hgqCGKKMIb
A7TlgFg28RQzJsDI71fauElk0kq1ChRboNn0CLhastBlBnRE/qjnQeXlQz3t
aE6Za48YN/gEkA9IoIU9/AXWVJBv+iCZxD2uL9TPqlOWa6S8a75r2EHoK1+t
J3oihTuILWMgkRc/FtOaMLG97LB30XOESt2bGUUBMaqoTDXs7GV/f/xXOQDU
LZyNOFfTzR04aelo8U8twOWYWtilZ+Wr+1avB/Fu44Nl6vdwjLsnpN0EQsO7
JTCGxbf641IYCEV1OXFDWQQo5fOO+pslFR3HZYxq7mRAc4kybUntZp2wGdRJ
ybYDkh9m04Aqli6DAXulrsJIkGcM9Wgz6R42HnevbYbILgJX6uMyErmWHnj3
pnVCBLmGBsAWMmQVJFiuJX92vSQw1Ba70137f3Hfv5yKVXd61KbQ2qttVtGc
r2fLUg5y4sMRotIXGnol27g7kCJtzDpNukJdKbDzmJT+81WPZqciHdm6a8jk
pO5ksl8fE8o2gi9josL/ftrKkugKhQprfWiCyZeDJKf0tBdixLC7f3TcmFfL
mZq5V+tU5RF793L2WDGspRt4GgEhExoKrUBx1uDGTMvzHn6xtOFU8wEh7ea2
vbWyToMETUvBxJiH1jJQDA71NAu794e6s5v39n/uLKKRUGkJeTpmwdp713Ha
hwRPSZTcvAJs5+JhPxKhge75UIrXZLlzkM5TbkonTUW3h1zRUafDOUNF4DZO
dr/jUDJfPqdoLj+LKtPpvp8dIbg+p04gkCBG84qSMc7AqGfb2unPVKpI/aLF
MKQz4HeN0gZaUd5SHJdaUSZL0+VEp1VzWn+ccWwuM+nTrj6BQFREIAumPUFr
KE/NWEoceNQLOZVYNTsUBl0wH5CdALqpJ3oBCEoWgnz03oT2ie+9uB0IEJ5E
99ad4ftOmNgXee2zUX0L0QMI0MDseOZ21tZ9NohcXQanf33wHlDJkjBsCIfD
8MSoo0vHOF8t5uDRH4fDhcC7GDNHXEyJVPt12RzUa3SKK+N5KUB4VEisduww
km9HO1Z3PqxI28pTApYfVjsI45AhzME+pkWLXmyT2YY8pb3v7Y2qeFniV7hU
7s209/yBEVzPgpRXPLLjnqd9i9wZzRpXCIu4y5tYL4HAmB2a14zoVL2SCUO+
PhMksdm9BFaCSFPMb6QKWEvunzDna8u4pzyrKMrVrSDpLTw9R/h+VSUj6lbk
SFZxVA38lDd2L7r0cqrTfJAlQ3VVfdo9/wyhCNJW2n+Shse8SXwzMBnRtLRQ
I1iNzB+mfUcKHFZJnA9ZjcWYVyH8lS4cszkLHWt5R0iqT6c7XTHoS+lrpdj4
NvIlzylSdOPDvEJfpQWCPvt6j9yfn1LNCThqUfPfbRlE/MQgKJmZFfDsPNnA
J16/2vN7BpTMXBsh6Ww/PobCiTklUcKqTQk1vRSMuniZxYORd+P9kc8mZmUX
WeGeWm1QP98Vjm6yJD084CXlLLAv/OlPSCw5Mhw16QIYr8GjNciCY2Su3Ihu
oimSSVmJDg1Vg/sM6iSMaEv7bb08Vlco37puMy3QtUHhNOsGNW/xuStEOueZ
xf7DPgPGe/qwYk6m9NL/V02vS8TFb4HuIN4YcRVinoVOwJngmShVoIETxxTe
tdiQQJwphaMjwUyzWaAelLWaKOblRd1Z+VXSKweXarR9WvdoXZghgRuyRvlU
ScCLMsrVCT4CtqDK1zHeG1JClYpCZoUtm0uDqollpBcL3bP6hG5XMpgXvg9B
bvltp+S4WOj+G645zZGUsJFNFGpxADAVzXL5S//VS7WCMC/ljRsLdpig7LLv
qD/yOiLfd9G4PWmCxuAHA8p2ntYqXf9dU6KsBfbx59xWZUKuGTgEn/za0jB5
OzEyGhGmEeK3MywewhTExmgPqWrQ1slosJzBO2RkJL/8/DifS6JveXElgoeF
XvYQaddy/vcJnioJm/SFhRj5afuXfZrpqs4BQ2xxrtEDLAL+qc11f/TD1U4/
mI31u0zRRA1tdcjvfyjxUmQO5L4cw6wQGjuf1vL85peLhAqAB7JJ4OH69/H4
cUZXhXnaNBo5nZ81kLGDmfl4pgQA5jIFo83JCCNFlwA7DRQC8AcsIZ72Gk8d
ol9kPSp89i5Ui04ZOSYHmbfa/f2ku7r8Th8vgf8LmQu5QFRj36Qjunhw+GkZ
8zxSOzMJWltr8tCI8AlMiWW4isoFFQMBOtowc8I0YU3riwldKLCLM+Ndpcb9
atxgNUdyMQKAXnES8oQ3jqEYZcPybSj/J85EmoJZLDOm1rlA6m+ztkmqD9dR
BeZ/95so5uZhEeSZqrkmiU8e8kF0kd2UQH0zkhPXIJlFHx+lCxLnuz4RPobn
D6I+FYw6FuVaO3PnigLNMkj9974BKqvfk+20ecAddha3z5mjrgTJmz2uWjvy
js2vekNEfifgG7Vik7Fgk5THkDp5ddyCDMHdeqFLc40FdiwPomQBdp10IRal
siETN3pniDPLufdjPkwLsZV6SqaixVGg32mX2TT0yLl80YuxYf6HoOEMgd3U
v8ADis0v0MoptJCIOeIO/2lDCiT+2a9BMowPJ3Pz4rN1t3ip2cHf26u/KZ8d
I72B+v9Exk+mME4afT89fFqNmCqNu7HJXPiBXaCEo/P80qxHMx0qZB/hwXrG
kjuFHUPyDUPpUZVC/yvXu+s2QK/p7G07mJKC/X8LBJLbQTN0TTJWHrKitY+e
L6D3D0dYeBNzyRnzOTn9y4WJ12/9rUFR89oMAJ2YboI6kb/Ju7gSkoxBrC9e
SqUK4dzSB9DuNQCat/t8dmZLwJ8LMpv/AqkD1DWxMZgOFwyGiVElWIalqMN/
lUois2ccBpR8moMs50KRId3BtHq5UKxSJKAQfgYrNkIdK/UqdMkgdMdrTz58
GigHZOm6rTw9o5G0avohq81aErIibO3D34EnrsjtM5kPcnFC6JdnL4plBnVd
GSFXTHF8XPYQaKiVn6lymDhmMPYpm6nHg2P716eX4bRgKKipvLHu523tL65D
21vlty6YvlcTfdWkwoX6vUJIigexELN9XXAkYHDrYMzKj8W7oX29SdTLKKgy
4ExlSsB0nx5653MuIPsVLdWaFald1P/5nnOJcEOgIeuhJg6z49obr5oJkhFc
0dfHUYdXxOE86irtbgQEBU1Lk6uyAOM54m3Mtm4fW25WwBeCQpSq8VY770mj
mYSFOra+EYIF/5Za28J8QdEPhsxqdhe3hy3qIoNzgNRQV7/bWm06+P0/UwCN
3N3ja9ial0QtRdyXOvCBnTyHESXldPirwlh4M5O2uis2KDli0Sj/chawOrMF
xkIcUW4ib6YKEnPfsx0Sbp5NlMhqWvk96wrm08rKfIIL3QyOyuqJweH89qr7
x6KsoMsO9Q+fHPzfzK2PRCVGRwN+iKYOQGEjRf3bu6GvZ+gmsOXhzFdaDUdi
1NMGIKv6fU0eVwVFR7IzPONiaRfeIx72flpPzzlQp+d3S1SQlkMLYLyMA/I4
WtQPHNstFoJgajwss3xDO9Uq3NiQQrdY058bucHErzEDrGxqv/qXdG1kwv0+
trRBaQ+k58mvt4dtAxnlTMkh9b9Q0BGp0s2V4uqlS/KnDJXefcYbxRlYebAc
sTwgBiXWA4/irzV/KryhBKiWVinbqswVb5EcMCvcaltkm+IkFCFxBQP17HFT
5rk/grMWTY4BPlUIsW+c8o3z

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NdOh/z3LGtaoyYmSC+C5BVVnr0UAb1ltTHwAhIFCaqEz6kGoYkY6ediorH+Pkty4P5IckEz08IGB28/SMfP9I/PHMhE9lbJVYr6R4FPCLMzhT91Lo735SBGekk4rkgoebNeUyj8aY48r+doq6izRITr0ceVBf5y4K5Q93CbDlDhY9IWU8HWRKms01EECvSlyhl5r6DrDKQpIJvLOC1oCW6Iw5ooE0PgmnqlRjlCA/eq50DOVFh8nEX0LrgouIHwLIb49XAqbF4d+Cr4M65PjgVAtMLgt+9cA8r+I11im49zZTKPeitNf0uLCwDkD3brIEVYZRCSSHpiiON/mRvOd/PU++27DpghkPhmK3L39ypIHM9Xp1Tfjlg4zl+JaOr5mo8pF8OlIyt2hTR4U6J9henMkZUx8WHJCdA3yzKzKi38yhMOWRNoN3yUKgn/tBfW5FNMwjKA6Pc9s8ur1LNdt/CAKKz7Uu3Gidg4sozbJw1My9u4dWdEYrFY5mDZZEQv9uIt9kesC3TSN04Bdrt19zIVyY84xDBDpvKuVUIDAMgrUHH3FDUtsaG4tJ5K8ZOiauDjOPT2B2MHZQ7TFBAQ5D7ITk7tHISdO9iMvES7DuMRkXPbVo0JdKD2fnyAWC9ueuVsvUieWJIl3emiOVhfNsz8SXeFrjfGk2Pggr+O0Mo0+BxXVNJCZkhJHS+/9MGjUd8/ApqZ9LWw0h15TBoxsK3xfK0Zdr1r+QUcRx3MCHvYj5kcDZ5Tmv6Ggjali1ucFIHYE2tIoTE1Tp39l/ef0Kp8s558QCifEES4Sp1WwxBFlYhJNrql1Tyzey9pe3sX1paz8OEPpQnXlVP6V/mrJeIOMKU0nw9VM+SzATRoUUUcF/9gIK9bvhbCAL4iAt3T3lpJaNnXYmMuziULvNSVp3BbTdf6/FsmY/pVSliH7tswFlrAg6QulvLsCcGpTkOCi8PzC9H50gVN2XaITANx4NuE/4fEw0Lm49pb+H1bWd6abTydbmTZ8rG7owk+0Bso+"
`endif
//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PS6gVqtLNXjvglAyJLEB/ss7yctcBgPf1Dpoij4yuOqc4WW0Bs9xHVxk8XZa
8Jqq2nkqD50VWeISN8a+NrM8lW4cZlBoYkW3LTfNvUyUnDf2tMsW850eIAc+
YfCwrsD9TxBPD9TgJCN6A93QsdzByyTWhnRjWKeVwMgqnNXwKbH/NToNkugR
eUC03fXOWV5GTgnB+zpxoJd2yWvU3/y88HC3iluMaPM8NK7WWBk0H0m53xbs
uK41DTVjiv4NjoE9YPdSPEPcpIUfcxCyJHfw/XOMAb7stnQagKA2yj2ayc/a
jfLo2zwoW/D8PKkegKVZXFR0IhtDnzPB3DTmqzz/DQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ebSGIv7sDcpnw549zmtN8IXqyV+bG/JbXWKI6j/6y7S37KyzIdrsPOFn+h1A
uD2zV97ZcRPN8AfKp3pnVsxqQStLZQRxLPy1bZghbTRk/q9j6TO/UMGJN/Ak
+wX0IJxm8XTfZkKvn7TMhyOHwzIVZHJmfG372NIkkifLa7vy04y2C3SpH+qd
+C0CGSisXIpQEBR83FiGRNiRbOks2TdB2p7upPA3WIHGAIcl4Xi+TVEszke8
SVKS7eJZuMd0PVwBNmx4uMlwpF1O/jIPGXpXJiCOFXdUNfzah91/Iw3XZxsb
tBguxUV12TwmZjm1gNB5R3tjuou4KHcb06hh/8BPxA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pQBnxjVzsXiMW2J0IczE2gGuj8mlox2LtLRGAejLSp1kn9RnaynqBm3oJqHg
WtNx/0vetHYEJc/v9zrAHXToPitCrIcENdYXCtb8MaalRy1bHGHg7Beh2lT+
5c/cnU3eekdT+B6R2lvpI85Yr3mAX2EJoyOGSk0hg5QvawuP4baiWGsqwf7q
kCTCdWFL5VOfR6b1Aa4U9Ru4lvglA2pEk+V8EeFH0bZs8zz6zej7TM65ovss
neyHklMAgGchxAULJDoa37aAEkUmJStbHT26Nm67FQyE14xt4lfe32pWrd1v
g+xlYOFGcJTyShLhVtAo88nwBC2i/sCZ7K5UY3Z0TA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VwyxBLPP8DPQtdB/cM7zLtSkUlgrDjsGExqVTCMCjII6qwYUTGlFFj1qQMfU
m+2Oin/j3YF0gMxFTKlB0EyINzkjK3zqbf368sSo9ct/3aFIXOMM9iRTkFS3
4PWhp1gENq2H91Yq+83cJSE4dmO/dwh785w7jW9BVCeajX8C8wEnrByx6ifS
lG4QqYWszQGKpiavJcFL2+2NwDiaIry1Mv/j7zdvmGzoivASNZ33apymvAw9
JWprjklFpjorSlgq69DE8gOA6hq+JJdh8xoBbkKcx7ijgPyM7Mry80fU9QDf
YGUbkv4PJRv1RAbpfik2fNG2r4XlVPEo7sdgrdpBfQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z1YfcUwOTtgKmJS2ddfUnBbXSC4Vfuqu4dpAg/PVvHS/fJ9pdGh3llGKyIzy
VEV3JO+QDxmzAqxJqV0s1vKdiJ40XJIFB1YVbQ5L4B8LL15ChrQQBfp14QyL
90pt9dM95RngWYycIASxUr+lKdMoPShmDsHuFNYodnEMYZ+JaTY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
r9RGjaZvYnm+rUwocuc77uF1NsYoUMZLAjIhkKgj9tPzZHoWUVQEoU1623G2
OBvTuXV6AWaln2R0QZrPwAeedTJ199K5mZfpIZI6Ymu3VOwoTLS/hzTtfc5y
Solq0wVpo+qHh3/+NYgk7GbMcqm5qTW2gDPHUE68fCnrkIBT1O+OpkapIjHI
Zt6oDtld5l1T3XhW+02DRrnUahr1v2PY02pLoiTnuq64ln+2r5xdV7e5gY+W
siOOFAFTJ64lRpPnseO8/qJOforz46YOXezp157bxP2RBocbNF4eQ07kcypw
gr6eX+pwTGXKhj6BgsF7c+DZBxse4ywHePDYFD4RjP8vHKvvpaFlfjqA9293
SxGd6+uN2OULaBqJY7lWdoZlJ2RUiA0j3z0RhaNq6KXsu4J8DiM4bWDO9I4O
WGMl+8oBRZfZQKAvVcpGTTOCqmmTwVEkZg6RI1SevDm0LoPgHfE1WznmQvlj
pfT5BIAuADHulrGLK8i99R3jSUz7oyVS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PmOFfZ0zz0gY9RiDUzDhaD56dxZ9yzTQ458NhW69eyvdkPuHrcNtXFM8yaQH
VKn/sshYSguE8UHsPJON4+3PDEt/ZfU3+Ihsa/X7Zwr9CMpCG6IXEACp5MrJ
1fUIpla4GzHpRLS7XhJk7LJxQtP2mplaJiWwy3iK8w4i1LDTATM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jyKJqSf1oYHL1QK3kkDGTsRYNr/Nyr1d52pYFxIdhYKbvz4/mwrC34g6cre+
8MYcwJjkA1udr2wuwU8StW3PHtAzQdVbNbLp28ns39cWXHRmDpd2P/0f5sw7
SP7AmbyzT5yCvr5RCi5PDAtXOtgTZh3y1uVwUG2QAzbBSvdf5tk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10512)
`pragma protect data_block
fPnaTXxiM5IkzDD8wIXnGkLOCvxuRSqdPyB6jKt++6x8pWwSVl4xHAmDaOdd
3qTU0Sd2O/5IFqux9N5mcwMJihhOjpNGLJh2O51LNHRK7jgLtlM+PVMW63Qk
owdR6cBfOfuJDpkuPPNu1FqM70sk/Ldaj3SJU07OIFpTAYhVYw2Ikx+1dtHG
I6UyS9wYV05O0zGuopS2rMSDG1YvH5UMM8WGJEgCHt0D9vVgQkSydhAg25J7
UpA2Vum4cy+dZWjHco2SLqsBbLz6450uuAY1VYb6gbhsCuEcEtGGqMiqE4wt
0VO3e4IXq/6xpU5KNQg2+CkNEfrkeHidOx1S7RXqkz6y6uhGPiGGiVSGyyLT
EFCn/BnSWMVBmKM5eqyX3OJbTYoPcenHmuHqRldJvRzeSA74hCo9P2IlKC5g
PDGtPRXCJiZcs8KnSaDfoe1Gp0uu2B9d4wHjHO/girXK3BQnbBH+fD1d6W5a
yEc0NFcY7UIp6MAjupmL9ffpvnjaYf/SAdzLNx5w+Mdb4mPiJ5TqDkGWbwiM
kSA/4QBQkxliX0zguLMFkPxgoIJ/XzwzA0ZWT29zRH8aGGOMJH72hyIZMXqA
PG3NYr5UsUQPbuP7BLS5qhtFpgBZNRUHeKXRdp9LpCviN9AEUpq1BVu2uRSt
sSztFgokw7QiNkpIJ8PxZVZ7tYGqZ1ABJZ7rZmzKMY8FZgqVSS+fCh3NuH32
dqDRR1x5wcftAAPHqLxrDNmaRRxOTq2w04fi4FWDG2IVAQWYmmTzfmlijZYs
nBOc8lm2MQ2OgUxGS9gegMIE4gWomhP/ukVL0phMUrBs1fqaY9xG51mCOo3J
EhVP2ZWGDxXGGd/bnkBLXefqmxN1fvA2JHTIrKTdEAlkpjfHyJHeL1iCjPAd
nc1dDFi0p+sFIWuVH7vjrr4hrW+/DIe6fy/sET12eEg0w8uRc8+nGgS5P3Hp
HDqEILHNVXlX9cXdxHXJVFK+BV47BW0F5y/zBUGJyhOqUg7D72oZH7OZb+pq
yt8Xi4Bkcl7KKDc76ieqFfPv+FuearQGQQaV6ouZ9Lde3f+NoQ4onvscjIl2
HMMCWVNCIwyKWLBehxk0VPLJ8Kwpbt4oS/czp9uk0PAxDzJl1QrSauSF9ZZj
r9kyF3Gu7/IS4yixnybgBNih4XgNniRjum9O3//vm4SWRhxcSmc8Z7Tlwyvw
L4UReNZLlbFjbu9ZGOWaWCqpx2S8K0kgn7ekn/i/9K9R/cSZOSOglSI0O79b
vT2fWwZURc3D09SLGzntOr+E9EmVoxZIS+aQSmvTvsYZSZ9lFgD9KTNRIs4N
E0PXymAldcNLRbL28dV8Z+avNN6q5foK/emS+VSptkuh/r5MBXkfIY02EH5/
86eUx3mPVfa6o167gQpnes+fMRR5nl6t/n4iz1hlr8vt5Luo+Beeocc2CQwU
RfPAuf2WlX7KbVzNakwclNIPDhTc67vl74fMSwMZjcyRnomNdjXT6sV/xLO4
rMH2EYr60WLyxdFHqECQ0KKp1TcisRLMRmhuSbFMYcuUsDjUDv8NnmgxMn2p
Fibowa099xTcfxW0OfLa5ZJbScSd5dLK66hTOwwFjk3AhdBPDMc6rDxptSrS
j9t2QC40pRgzjFY30b1BgaR5UbedGUKxqmcROx1hh3eJTmdNZLZMBUoem+et
jqaOUd27+29JTNTrEYJdn7hpKUy7QhqFUIcaaCIPZcardBHRZg4D+d+m3iHJ
xHPr5Nnmy+5Ov0wOXnHoEJnY+dNlVCEKCYdEBQwSKAE5BsQYezaHe2dSnPzM
7vgrIbjym8K1cyV36JZ+bjsw3TLDZ+A+iD24V1PeyQx6mqNbNPwDm0zNRQpe
dIusG4p2+ZWmv2EYdjdowpIISv2dNa4s0FSs6ONmxgkZmlLQFDZ6YKJyHewa
rH+66W9YtOaE/iOJfyfosWHLpy1ttp8oqhPjlCVf2j6JDk6CzaU9bhSmj9mZ
ecLTSpEgUUx90K9bN1m9nOMX9cjZMT4OyKHYujK7Ryk9Zbj7dinLF7IIHo4s
m3n4kA72anC22eqf3+8Nt32YluZCtLBe6r+fkgCfPLKcIG/4unk2XJtJP8BR
ysQ21T0TTLTrEf0c9jMMWtzWs7kujkp2susTwC2ogubByK0iTl6DsqfDJP/G
9OzBihcR4lFVyW3LAFJyWRhhnFmaQcF6xk1LCp1+gveDoGR0rOBmPOLswvaX
r8lnFkpbXb9zn5trWZKQD/pdH2OSClpp148inZfP2sggpvylB/76nivilk0H
84uExG92emRsbIMrsDotfzxPNiYjzy4BhVgRcpDwmyZxAj3xHUdSSqIJG7yh
fHb+Fyy3d64Xx/NQZ2VSTSS/XJbh8+hRkzBt+xjy5U2WCKiOLCIZhwIuVcrD
EVuZi10HurRf00J8dFIA75aFqVps08k3C6n2dQflT2EDs7XEMVMHFBUVq9GU
gIvNuR6YWhHDcQqIWLE5zjr22JbghZIU1/vmHaWBz0uJkx4TUO1pSw0V2KGl
mly+J72cegX0N28IGCUIU2mDMRY5sVu85+pTkjsLZLFM4ZcMxRlkmJ2VDZ2b
YgPt9ISTUNWxzEaOOAlwuCfRK/dmAw6+R0R9Aa0Kfo8ycPlhI4qSWZ+kwKbk
hkMQIA6CaQCnBD1u/Oi1YEDs0Nqxo/+UWuLKggBpa6xwtk+N/PhpHhq3lh2a
FC31d6C3OWNX13zJUG0uJS8nNozJuhx3r7nmSozMEp+cj9YTnB5z4+1S44nu
QjAs7VMJxPGD6vW07o3hRIqYmHFxnaXtoDoZxLy18xyExeCYILTNt+/HsiF/
fF4GGoNTWGbWlowTkn1TXq/uXSA70UD7TaU9cN3cobkBw9NJbEe4xFZOo7J1
lzkawlGaFO21Zo8+cfdoquYEvcDKN7OigpfXQ+HCkig+HRu0MPXEOrOvHbEE
Zv8cRj98NqLpegCdEE9zJ5BFKyT552xgp31nmDbl/e3OnFlTteLBDk/l7TDQ
6y5xLZzRIDoAB0TcV7eeOzX4L1FtrvqUGMRckgBK9++gXVkRhbOFHDuFJBgL
c6q3Cd3OGFNZeHKOdtr6j8Oj1noJ+CmZzTZdIM5FkpI5fMcystvVWoXlJ9ay
qcoY83VXdRrjsh5/FmNVQBgQA74ag2SOBOV6K4imGdpKSntiQ0UNiM8OtJre
GDWrtgGKajf0lyqlLvWSQAaRkcO2e7MlpyUUSlrmfct0N3f9JpBV/1XG9RBh
Jcru/IzO0CpvCZOH3JmG/LPjGETJZXZM5x3NTSJLQSt61ESfMGljPOhVpDr7
xB/B3AoupjTCQb8VfjooZMYI5040MTISp2tAvbhIc17UwnEHKDl086bmfDey
nWLhEO/U7kNVTzTud3Wh5bvqdS4F0ppiaYCyRKUeIaFOAnuVomWCKcAXFYzO
vBlLT6cJD1/HJcKH4/8WsGGAHtQec5RAGA2ZAkFtHjCj7R/Vdgc+vXKdTwAU
k243Gu5+D6s813xyH0EYTAvc+J04zQmmJRvIibbLGv0msxG+2bpokADsvBpY
1CNxpVprgD8a8fzaOMkRbmqVF/552iD5R4fpTupTMkRugQ/wen8/tg/Jhcbu
48JqVpZwAu6HX85Ogqn5uvydRv4T6S2XA1fPY7iskuR1cTdEn6emGrR2Wh2f
Lv5B2EV9YIguNSId2bgyMPjqzhW7cdW4bUHj2r6LwHs7AmrNrWrzOJTmoxVl
hq+4G0KLEBu7oauQ2CNdKr39NfxL1BaG8v0vAtzkhR6OUhwjSLPXFGlctD+S
DcGcI6i+8IOFwD06d8zieEcD+VTRTLxpxYHDyvgso8dFO2dkf0uJ4MTzXkZq
n6AWa4O+CgMjcPvG0jTiuY3ZOuf7fnZlGfDyQjYEAieWBsWYsFhiaTiIUlGg
ieOIgiteXbeJLjg5qrBvLiwFibNsTkuOpNwPUToavD1oLPaQFRZrdg1/Rtpz
SrbQwnZZ/TuGoXUV3zPESlD9fTk3G2xIgVQS9MjwZHTHOkUFfRooSsK038Xm
ojlPDM4D4Hc/BSJR9ChCGKFlJmpM2ODpxs9uGYeaxLVde/VGyh7diAIZuNRe
cYkJBgueKYE84w9dQexnveG+Wj3ca7jkyO2d8utM53H2eMuQBMTuM7CpYFs+
MLTSJnFBQnb/MDn0VFWSkQ/r1t1lufwcjdMC6aMGw6IZ2gk6Bd9IlElAW/+2
I2KH5rq+AUNe6je/OAPQKdBvSrGzf7q257yeC1NqdFdN/LAMCvWoc3Z1SCYZ
9J7Sh5v1BudlDWEDFTXVckLRL1Yb8mMuACLxgFNn1RJdlLP46KQmDt53/Mcm
YYM2l+Ys+mr+ac3oPoaQwfwCDSh8+HTi/i3yXSYxqMUAw1+WHEHtO73/zp9E
HuZ717ey1WR4JoE80p81W9PXqhm37rns4FEOY760K0Kjb5pOlAiucqkI/cOM
f958xDRZ0LdgKnPwbyXLAzmF2c8UoZ3qYxX1Q2dSHvT+Hr+NI028CmN83imi
vRelMNDFzJ2IUHwQmPJXI1ca5Yqh3MJxAcGBpp4ax5A0La+j7/KsIJ7ndXrP
6u4DfZq67PZar8w5HAHpxtDlAG1Qa6CakmM196O3c0mdffFnDjNtHnX+D+HK
BqrpWHX1nAu6t6S11zlZjZvvKoGZ+FGtl2HRtJZ+Zuztq04GaFzCvunSUfwz
kiveHB+ykM3AHRFwhNhNhHBVVDe/EAaCjPbjRiodRR/GWOu+RRenE0+Ut4mw
SrnLMupibqLxW09eeDWh/gIrTEkYdSSyskDfRhyZDt8hXvZzJ4b/KG/LTgRy
yQyPRUwDJGE8IAYaphrYP+wzpAhIiUALrQfurdE0QoGSZd/aFxUjG0eVWl7Y
zMinJN/gilRfzlJ2DpTcf7P3dOAleqUCaqc44YR76Ox7P6ZbhHl3QztlTTGZ
pXuhBIhacu8RWe+wznAh+/YFDZu+48PDJprHBDQVP0duJbY2nUOhCNsac3dX
g2mqX6GPbuTUszoWKfR1OESdwpSui1HvkdptAlgX0LuoFIeCZzKEVuNQ3pFO
qH6QwXO1x0ikGACCPb07HMi30Kzk8+aISZNYhobWZuBy155XKbmDksuvQliJ
bo95Oc3pnmeK7b/mDE6hNiBvqcRbfGEL34ZMpTb9ETmge4bYJzIptxKVfRKx
YkMgkRjd+ejgRU2I+iW/0dSr40S1xz/MfylOgeg3/DBE62SHnpxMYjSG2vhM
buNu+Mi5rDRWlM/MCEOuEvrHoE2qvFNmolp8CMKOU/cuLYfJw25UL6qYOyA2
jwcYCX5QW7w0zVQ+xavhafwWV8yzpk9d9Oto7jZnzhm3diRwWRTnNLTOEwFY
QFkAepuqj76w4LA7Tlq1Kc8eUe6V9oRghAjTics8Yzc8ieWg+7VR9LhYAa2i
GBCiIYdIL1ABkoA5X/WWxHMq2m3lrhxeWZY8Ag1XXIbVgdC21vODslMWWz3U
rPYQpE/nOLqsm/ApnSp19vCWL2UBPtHgRGswH0IgPn4WbpvY1CgiMs6l4gq/
PqsNXV8tEd5Fqcw1xLdtaaqx9Wt+UCURtydI/spGrc7omaPFbs9RSodwmHKM
3FoIiQRM4BK07xeovDJciQ38NB9YxyaBp6CHeoabXatNwislgyS3qs4f+F0F
tnMt6ho7NzuPPuFoUv8uEYCsI/qaA7+Fx7M3JRJSWN9xrayJvF4TzDngoAA+
wObcnEmWAqRphTREaREpawzzWaXPvDQpJzPr9Qqb+bQyJu8JFOAfg9Cwm6h9
PYwbrCbAOsPVecaLKTb0+WrGEn929FPvHt1ksEdydIJO/R34VMgJavRcBjAa
rBP5JQ7DkCJkUQiZdacYpI863E7YGDbfs60SXhdZzsGeFR8WzzaiS4lrzFTI
JvgR03iTggoDMcc46ovFvEusrLNxH7wJcjLYy1FFZSyqGzCMIXdTwcwjHAU4
2UdFcKBkgS8v1LRLkijQY0eUUvRzT8RZPZ8l+ukfJZSu94ymgS2sjw/MJcaM
Jx8w4wBa0292sP9eMHW9L/nQdAqkyDyMt5PI84Ao9bQbFDF79CUFFue/RVa8
a0KT6VpQH9aHRjZ/UMNXuOl9VtUdVHnP2C4iJjyFCJWoMzgcYhYMlTrU+12k
4+NvUzfNiEGQa05dQkmEe8sIL9r6YIdVnmFd+kQhXopd3H7Uc57hORYUaTHx
bnoNJop2LgMBY8xRj3hn7hfR3p7bi0cUnGEIo6KI5mSWq7TI6QN9t55OOku6
bK3FN/9uUwYHBGF8NLlQ4X9DW2ap+lf+IlgMDDtjZ94cCrfy04CEfGCOLt9X
GygNqpkHaA8VzjN2sFlVq00OyX3n8MOX+AhiqiMWo+kqcoUJymzZKrk2nza3
Dt9ckou36qrel3bpymdog+z7sz2dqKHCFK9Q3k+866XOWNP06YNEZnItJAuA
uGLw4RFCCF+h/CnpWqM0DgvkKBuQPqxkHBAP+yKTDwNT5cCzlyNikovuZZqy
IRIVLfFW3TfFKgYh1qWd5z5BM2hGkjO49exQ4pM3DdV4dwiB0erX2hHc8NY7
3kDsGUXivBnLeQL+ELshDJR36H6nKZgLgxfNRuAPIiLpy41Ky6/UyxfXUnI3
XLNtE1zobay49Tpb5rWcREhgdfG2iQd+Ef29B9/aECArIMMcIDu0CH8sAwVf
MvaW9hF/k6YOa+S7f2UA/jY38NW/jcxt3GIq0z3XHk12tCkH+UsIMKI0Z2UP
231VaXNT6ZklhuG9Rr1eGvFOrhdzaYUg4NFDS1YNxGBZQ8mUMpkod6UQG9GA
1t7wbJ6l9ifBtDbAp2i5E6yaLDaEN+sCY+AeRwkoBjf3qoo8BGUX0e2/vrQS
1PD2Zqvx72MrZNTdZUwiUJdvZ59oqX1/NXExLlVwHvNYCk6z2YfVGM9wLvA3
yM7+nP82ji6Tl9zda5vjsfzasVM9X/OqZZadc0nghPV+xwY+rn5YX9HJMYcE
S3LnnabFHBfAK4mOXaPeXIbgu3jE4kQgzEpAveZGZ/26P8mS7TLKc2yGmE3g
9crFsAYMAS3idwI/Qw45Od7D09A5fveJQe0SsH0DB2rvmtjJzlczlnx+oXDC
aNPqBhKQW7anGgCnjMxKle18arUCmMgxTgD5nfkOnxeVJZcji6cMo27sfxCf
6K0NQMoKgdOeVoUjk3vArfnDYF3I59W8JWShFQp25fIbxpSH5s3ikTfWgC1r
o1SuqCOGM3vu96MtKs2D0F89ka/t/9yBszJnxT/zNB/WFZx4c38tWDoLeBg9
lyp/p1KbQ4ZE+hqljYjOdeDiO8H9aapdqnI+TY+dQ4loqfWDhkxAiOqYO30k
ux3TrhWGeOttus93wnhrJ7cnxi4V2HsB3lznlCqWt1zd0dZo6FY6dBX0Dnl8
/iadpVbtn//unQUxRxY92M/1sfANFtIgky0doTSrM1pmEWs8Fxf/i6N+eAUq
P86wqPvPZtjicW94rUHoPCcD7EsQaYmS7F3Wf/f6RiSZ0N75SUNBIsxEzHIZ
jZPpZ0HyERa7eFCz6DUzbjtDzWXIyxj69ad7Vuo7Bc7VbcBwfpAjXOYIIqpr
OYMfL1v36DNqKB6bnlJsT/PvQKEi9dafxrAHUTntCid/mVAqwW1cK0P9QmWp
gPWnBfc0a0xcqZJDxC8/1qPL0mmkM0QEjDGhhStt8cmoq+opdbWYhiug4t6I
ecJVI5ZGbDoSWSvZjOkfLsaaESg6Vd1q5el+oYyuxTPD9KCwtz1LoDSZBL93
1IzddrW+l89FUWq74GHmMSrYx1o65kRnJSiVPOYQHhbzNZnPUVatGjAUdFjj
yMCbtb7kjHgfDt5uoewgo0+0NIOkhxUFeb5BqhNKRPPLmudPYYIznkz1FTTM
TbuUABgg+dRjz/lvh8oC7PKBnrU+NJzxhwwX2cWCCjHeHxE07s5ErOgQQWI9
7M0JCrFDNJZA5QuwRzXdsFFLBPAB8WKW2AqoqLVk2ViP99+UX5md/Knv5S6p
zpfjGPBTfOneHPLRpqHt0Mj2nHEV6jZpH2pW4ubBvrDrW9i04PSmn9JkRP6A
UO8d/zpGX+hcHWrJw7+cyrwXamMJtEMYZ8EI5n2aX5Fnw92PeWUS6O6fWS2C
/m701Wjc4x5pNARk91NyVXDuVXKbrwAEjeEY4cnZUVGh48dsyq/uTIcXTjtA
erhjriUV7TWzayQcfJzjeAR1TbvC65c7+OXoAtS7zLqiXkAikkDaqdGio4S6
cNqznNbBFE0s9i65kdxJez9ygzB/wS6YhneLJkdKzAa0DqrQBHy9evvVimzw
ceIEeO94sO2mBJyZTkjXzgXULvnyF83Wr2Hun+QxNhHvXeTcdWeH+KT3ost6
a7HbjsHEB2MXbTE+uctIrEU1jaHW/U6s7z9iY5wzMUT87ozE4FGPEDAeXBqP
4Nsmzh1CFIoZEu1LJ3DSaHFOsLpJCdA8GnaLYdmWUg+o0B1p+URGHgK8Pk7A
F/5FQPIueVj447Ps5XgsIwlRAcEM9lxcdWKFA07IOq3jRyhMLitaYmjI92Es
Yneqawdjxr5LzZBOthZL6yil7wO+yI7E4uhHyWg+4YeVlhvU667GfiD9Rwot
fR36Jh7vqNrQwk2VWC+PEfpK6WscwyfRsvEOu7L/SqrKZr9P/rjC4kIYnrgQ
Z/ZDgL+uOgctU33x8yhJlupRu1fBoyvn2xP7rAZgE4usXDj2TNAbl0P1c914
1iWl2uq0zMT2PdSTkpocwHC7UDKtNRS7WrZrHGbhoJiLf3AlLPCfKsPSpTma
knv4C5GsCTYTFVofuLafLsRxERP1ySNYz2ZQHJ2Z8cVbwqTjHVZdAr0PfB+c
Dpzq01/9q4sCyXvqAghlyR198eMismbsl2YaT1GG26JMTXqZZMREZOfkiBqx
ErMRaZWbl6wpSMVMG9wHBbA1cuySo7NRhUiNzO3gslyzSiKLLFv6yn/hQOHN
Lesg6nDxav5/hgCJDB3k0lo7GNdLDGSm1KOs51nlJkbwp6T/9HkICTXdPdNE
DPgk4itpPBg2bUrhiRg1STxl0twMV8zvUjpTnN9bXBBFZQlagJbD1JtpEuV9
+fGIiIIB8+xCDiYr79kZMkADg02caYMPEs/v4Pxp1SV5tId2odfb71991G9+
pJdSIsnZsyK0zqgt/T/DiQBqrbqkTzEnZ83qGdwHVa44VW4VkUqsSLB+mOpt
IEjyBrH2PrqPIZ6ltUWXzg+dde1N1gE8WPW9r1uyth/K4kIY6j1jrNjPW4a5
xtyt0xry8DgDlkXv0iGMqZgWdbY42tZUrG1L989YnJphm/N9E54tKyEQ9cvg
vONuRa9FTWXZWC0yH/fxb5MMqXLbT5+lDpsV/m0DlPMMfV78k0auN2vsDjvP
v91hWa7vO5h+k5hjziIGJp0t0d4yO2u+hyFBot5zC3Ea2cMcQJog+Akkdoev
YsBMxdGfSXidm1pe2uLjIwDpli/H+2XziSRnVbwaNhMC4eK3tVc8ZCbElsCn
vUThuzZ6PdWHgIv0WtzEWW334OXkm+YsFpKlQO+3R+BU883WanCJE82xbl5h
fSWoRNTg2V5xrQE9GOF+vDB6dSEbjT82aw43JAMhgQw8JJIcn5wLxGJ1J8vL
DMNdxcRWPesx93eM0M2jFBF7fxBctpVeVRbRH1VBR5qj4Owznn622CEenlwB
hM/6k2jEI6N6eqHdw8phq0N5FF1nhnPyW+AnWyb2VgVY//48a1g+rDcedZOc
SKPphrsbUIbkJHmLluT/oTgVF3D4U/RWSd1JrZEkzF7mIeuSBEr0LEAf/qPl
vPCO5wp8gLVwum84Uaw42RoLCmCz1TFrGkDHD+Pg6RVbOGUPjA4YbKjs3Y9S
Vz/T8OG1p5ZooCrwR4DfuRUV0fq/D9jKTG1gB2fZgIKgLgq6DRbkiZ7vlIQV
1ArmASJzVKCbAD03k/P76cO3Z6AfHZm0dussOz2+9yTCaK0be1bX7tICXEpW
czEOjr3+65yZk9xREnERaQx+QF5BzknB3AjBbgNW0KyLTXmYr7iQLMUXrIjl
xlyk/XUWv4X2opT2UvyD1W/KkKL5jXaYUQye754Gs95SAQmw/X8YlnorqDXU
Novi117AxHuebBkcYG3ez7iMKySlxZvvxu0Z45uxt83E1JB4eFbMyiQCmDzF
9CfhTawmC7ZBGaagIRmMIYaM2G9NNJFZ2Os/BHsGm3wdVFNTle3bmaK1L2sY
EvDtCo7Ky8U2vLbMIQnjwsnB1JUmL9WAUhCGvZtPyuED5tcYvQsg/q76NMDl
fW3+zK1YU0XsdYq1UfYTIw7vWhlEqiKyrfvUmkwOG41XX7ndTgLsT+F1st+R
CbzCkXu5qZ8nmWxx3MIIp9Ks+8l4x7p1xlJS+PWymp7WSn0Xq97m238tXNH8
rpJjrwj6Of++vpUu9W08a4tWzsrAxerQtR5ifhwDhzKbDP+jwC7IWR9dAk4M
UsUpVv6AItfBJEFAwV4MqE+AiXRt+r6LI1Kz3l3oksdiw5ZM0FOZbwcfiN//
ukmLm5nbJyELa+Zr/YK+wOuogCDXu1PkJLeRdbGyETbhCcDn+ArHmz4FuUSE
7GURLlJytbTFFqedfkAI53LYSfDK+xZwNFOU8OlUX05D3R7vufEMQSFkTq+T
HqR/m4xFmj0IEww0WWaiT5yLJCS0jwkT4JPEf0txf4FSdPfFAEC/pAAIrnCT
xZicxpvGBq92vIymBIgwi76ogjDIPOaf2AdMZnEiw+1dIi1y9rAPi5az0N5E
aj9EjSGSISS8hgcNmt1LWRPMpsf0fjum39JBIgrIGQOPDYUw5PSewBYOI1Fl
LcllpcQfyH6+ImI0obaDl1DNjhFigAl9aW6F83mkg62jRTOiYMihNEXmIvvJ
9KyZBd6OrANvEg5A0mrICkCeDyR3jp7w/5yzGHeTdZ667PZtk53dIQqMEboe
ACjI1qRAdvlvdoYl+SW92/RUIb0cAc8vNu8wj5cb+FnUbylOp18o1sncvQdf
g6WpEcE5olsV5VO8DJqowh8ElrHU1+iDShcn+Jj8OgcVSx8SxJpIKVBN4FVc
xGYnrV9v300HXOBDMvgbRD+Wm8Yux2gQmon1agVbWs3MRSAQSfEjMcPRPGhO
AUWFQKw84UJKaP5kEAW9zpKnGsyyNCek0Tt3yki9UlzUNFr1WUvrgmB/oCxA
k6wHaIVueR2w27C/W4KYjbdjzprst4zHk6LYPQlZCGKaEV/8VFSSYnqsnmi7
Qf5gFx0BZkMIVBhwn8oKjwnor6GenLn+1gvYDDhWhnEl21DnKejZvDkz7rKJ
vAzneihNPQtpLvxMgsKo8iDM0H69/vd+Lyi0ypzbJv3DUB6KEcyngfcLPKo8
aFZML+tSlPLYmDHgMvCGfY2H+8TjFbhmO1AiIb/vmt9hCyXgc/q7QhZeT5wv
qIRNo5nMyMUdmfYaYfRuStIywnf4qi1B45e6PRHmAbO3LqgIlJgi7wZRIT/z
4yxdP+SBSwXM+MPh5xR5mW7v4nfeGQOjYDQwL7bOzIEeO+x6CnwjDjNvFHYg
6SVrFNJ+aZZF04sMWXHLTlsii1uHoYTG/DpBTAYfYKmssvnUnqoamQtekGt6
WnBQvPTE/YHrD0A7bJqivvZTmOIcIMQ8cJCda+MdIVNfJWuDCp3H6pugnMLD
awmNoN7EhORBCOZJO2tpP4TC9za+4A5LA54mUTnJkho2DwbQ9mGNzId2a1lu
yQmccUzPl14eZwTDJS96/eAp02YIeDhfKxXK/oV+dM/IvxFc40beyoO39e2H
tQyFURhKT9KbkOgOsPqZqYI3x88s0Bh++fK5+pj8Qhn2aPq+HcvN3BmReDb9
OhgFDRL8PilkRNM4J9nyr5LdgSqzEMbWx3VbBBmLP5qsaGRsDzjSzpc+zAce
z3GBxCSsOS9BlVioUCU5J29TxFTdPxD1gFPlh29rVxfHAvp2Uuixk9TQydEc
aSUShIaV1ZHljy6qEsraAS+ACn5GtYUV9zz/3/7HHUoRxptl+QLGl92ZOqXI
PI32L1g9yp1Yu+/YRtZIOaHOXE45R+aFUn3wdQq8w67q0bbjX+Z8iLZNUnl0
g46vCAx+T2/Q3diybPmkQEBj330IipoT3NzLHk5nNNNRnfjaHw5pEx/Dubwl
xIgcabnm3s/5nQ/B/nk/1tHMtIWDKZNlVoxPS2SuzYAZbl79ZROvU2XMs8+c
DbdrLoCXCe5q455YQU5eYpDFJ+NQPkc0nV7ctkWcimQEtfSU0T8uqJkAv4se
qbUZeDksTZCRg8dBKEPP8Sc434Khf9VFD4DG4+Uxa2L2LOPkH52JjDcm4Zl5
EV1MJ/DSxKO7umUMlCfgRoSY6wumS9YtRiQMaWgvoDBa9jZizbhvP9MC+TII
oZTB0QMSzl+r7jysMOGvrNBctK1yHydE8nIb/8Hykn2dgzCyaQivQqLNojY8
MYrP7W6k3rkLuBk2+BxOOFNIRfOD2DfkEOjBH5t2N42xTLet8jeXDS44A830
jIFLkPlcOLde+f/6xuYrJWU8BnaH08BOzx8aPrDPxG8O9YPNUHXid50MWtqa
jZDo5iSmXyzLLgew98ZSYDY7IxZ1gTqc0NZG81vYMxRrujk8+RQXKAWP0dDQ
VE5z9fVFAGE/ScTPB5ZTIOFisc63G4oqZoc+ra82rBdf8QJGAoPbpnsZwrGJ
Ui6tDA3JEbkwNf1LJQ8weGYo+dwXrNXkoo8KSyKTdte+wT475D1zceKP5XIL
XsmifljUPa9pqAR0Y8ygqWgZqp7D7u6SjoxTwt6a36dRnLpWNFX3r83K/haZ
fG6OSAUjv72Yo+6aFq6+h01CEgyHk0jcGXJQOJ/KSgYePSoxKFaz0BWgFzyL
P0mtSjQ5DZ+3E6LAPsWgBPIfFZ9+tkIwsF82HU6GDXDSEwuyff9+sLsg1UbI
U1tDY68hq9WmqUESPT90CJ+JjohuNgCHAklKHVx+JQxF+t8W+1rqgXxcBP1Q
RrygMYFvNlDZsK8+e8oPoTQ8nkV1fMpqJy1lbEJjHyRObPQaaQMVwUDLcJhp
foIs1/F/J1trm/6jlNpd/rMnvGsEKuhEutYovp1iZK4zSbTeYTtsMIpq9Mh/
x6EsFmnf7WeTKP3SHc39JjuUJrPIEpwFNVzKwTVHBPdi17Eb0hnjf4x17k5b
DonVe4K7lgBkfz5BDiLQqxqNZz5+x4wsB3ZwByJ2dGAYimTE8lAO2CRiTlqZ
HmuApg70I3pNkbmfAWwcIs9UMl0eLG4Lcoo7kTvLlYjKuRWdaUdCY4huUjwa
mep8YrF27XEGDORJb8HXEfEm3GAtGtbrKxHv5CsJeJgCQHCrItRug1nU693j
SAYlaWf6zNMw60N2zdiKTiDge9H7alkEaYY9JZ3VYbn9bIzG/aToxqV/0EE8
ngmvSngjvA8jrCQ/0VwHe0CjMz6yyXN3oXDBI189XP6QurZ/SQ8Zl0Rv6tSr
ydzgE0RXph02AGg4Lxg0W8DUSYf0k+UqKnDmH9FtNCAzepXYYNhMDG3nMH9I
Ag8BbLo/UFWNqTKmi67ixFVzLRYa2PJ1lJjhIwZshkmk1LXdEgie9MHn/5sm
HSw71XL2YnoKT3YxtjejjF7erkkkSqaY85/lzHfiKoqLLo49bwRcZFphQhY2
RWJkSqrOWvv21lnBQCgg6DBAeiW2yHJA1FnFEp/IStarxm+9Dvx5cmfpCgcj
PT4XVXDE2/TiyCptcYP5/6QplMdKyIIkVIFJ2KOz45XnYI3sm7iruabgsq2O
0LbGAKv8Kpn4usX0/fLSQFcrvIfTGBfM5bl9PrXq+ZphWSVuGrc3HpVBsvjm
sAKXtwCnLuRgEgfLtMc3aI1twSHEEqWUyXaGPFZQF+h2nHuqFk97gxOQhTpq
I1AwbRGuO9gW+1pqD8lVFnZsFCqWm9TpK0f5jdNBeqILR2mkprB1rmNCxhm2
1VTsHiMBJ+oQCHsZeEurpr9ibVrxTW7tUvH4bRmVjqCfEnc8NEfyG36My7Bm
EP/qCk1D9tZk2jelLeM1njD8Sj4P5WpWu2IG

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "1YFekphAtdNWmCiTRP2OoOj4dXM8nCSJWFcg8FK2oInJHC/kg/p2pkkaTmZrbUbXdcmJjcaOi7c95LpfF/xNlVlYggo9nClSlgHbHcwLYvg36JX26Fc1LGINgbtm5C200nd63mYO2zRr2wKTnRHPd10nPRAsfX4c3iGu/rkzRZ4YQDUPANGCStrM1MYmGdcX+LN+qxz4+HkwclAC+iwjet8kI49aHK4n58/g2EAoe750GiZ25zPlOmhVXexEtMwFQOzJcBSzmMvLiHgM2rm2XAJL4Ash6xdrd/VDDVow/Rx97WGD78VoLil+/fXtF/sVZ058Q5pWl/OeRNz+kMlN7pMuLW1FHD+Ds9Y9ZMjcHjqPs59x2HIRGQtPvLSLuMOnj9E0zMC81ZK+p6wgkeszHScPRmJSBUervGkSCeSaTUy0w6qiwZfukVv6rOdtUVrmqaYdrXo7kAclT2Tc0OdCFNazJh9SEt01asd7nRO5+hkFwEvWRZnko5yGy6hAF3c4+QtML+15TVApm/ejy/Vx7cZecgtPaf7FcmGT0MvOxP6yjsw3CqabCKuy5cWgOL9K3Zb2PIsoGWZrbPbXD8xlCBJ/Cdm/7rvhEl1f22tWWVt5WnMZ5dzRaeNUzs0yGVHg/b+/zXO/1Bljop2Azkafwu53UiSCjjFs6GLwrqEDu0QoveBotzK30U7UJ3e6zObu4qyckgKe3mfdQNzHzkxjPEy62DKx9tPaP8Hn1ZuIzNcyu49fbNyhHgvHI+QXxrvLSZKSDeDci9OpFTgwzdbuXIaT+3e+WeIgw4kjpatBLgHQpOV7ku+EV34WWviogXUgkv5lqFxBQ8RQ6q/DiIQ9Ye7JeLnbV32Zr4Jm/b83rq+l/PVhVEcoZ0jjr339biaVGndIcKqV+CIAKq9yzryKk300IAagccokhUu5OWzRqFd7YcwVNihDcYLI81S35gkO3fzk+J9OFqbYHgPLnMWHvXVikHlODeBUi11kB+julIFGfJQNd1QPjKP5JQozJhwe"
`endif
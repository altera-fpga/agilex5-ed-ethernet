//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K6J1MFrKrf1RhCTj7C9/TU3MYDl+T3bibOf+ehdeIGp5wBjX+NR8FCfR5KPL
LUaVFmrNOw0vV57SHPgFcTnhLniaAhJ+Q2e+kCjxdOxiY2YgW9mJlBMwHSXy
uwh2eKMAB+KJf9naRM3AUGKED6AMs072Y/5DaB7xY6u7t9jeDkEqDCgUN0S/
awdX7XWZDW9QAE+z6XpJ0uE+h57U8fl63BeaEQ6H9SyxFIZLGL3FxB+oDtoi
XxMntamigmIKZvPeIwLkBllq4Rb5MWFXlJ4qTuWm8MR8R/oEoNETc8F2QAWp
oV2pVdltZK48m9ot7p34d4ps1ndHZc5Zrp5l44TYCg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TcHV6Inldtcwlw1R4HpQGJL9Q889QEurEppKgSiZ9KUXSSiqqsS4GNw6FP0T
6Es8Sy8uA0kEnTm8fhmGVyXv/03jl4Oqq0hNFYQ0nm2G/e4fZhVrUyaDoWXT
VAB/BrIzDzFsbjxo1QtNLEshZuw8UKynE7V2AP2mrIArO6pAzX8Y05ATucCr
Ue28H07NpKoZVgGEyemC7NmQm8RCZNMu09FP2ricZBNgUZILvdPON9YUYtCz
iHXwuQQcKFIr65oahS3B4ou5RskAF22ZWrm5qM2duIg2rw6Pwlzg5WtK9CRr
Vm4XHdMOJoaiHssEOYJezBaRs3I39qDT9Pocx9grig==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
brTZ3bLGIFBqL3YZLUKTtixf5+IqZK/E+E645c1iG5HlXIXqukz+uE8iFZxy
4wvlAiCG3gXEk2JiGU1t1GfTLlr0x4BUKxm33HGkswqNVJ5Zk/gk8VeS0IK3
v/hy20ITIAi6RpGx3uXTqO5hXEoO+wy2qRGKXUfMtTwVzZj9ehzJ0WoESvdo
L2oOkjBqXK73PSXYsL98SC5/P19dPZOfzP3ULQa06fScWhO9Zt843vitga+x
a7sYma6itjWWQfSj47I25mRgImKazD381EGzWrwvbfgXW1AhO9UqVbVVeLt0
w3EhnPYidrSw0Wi3pZophtGnPhc7fQABT0o8NKAs8Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CX+MTCmfwoR1v4ndViviSxU1UuY1L4qShn88pEO5ln+uCWflYgyadKxAx59f
Z/sgbdCWPJ62OZI/TPZVQ5pxizdZQI6GEKUGCZdDc9mJvbXtUl/7YK73+oV3
ynK2t1N+AGVJJEY/fsT1GHBw/JpGa1Q40tYwYeX/ohmazLlnwVi5ZEaS7xAp
vtxUJfpI5CrIeGiNHIIHg0/oiFEK4APd8YsCQ7N07No9mTiPCyQSWC+XDSSu
+6im1JiTES9U+++sjLZvlajQNvQfNMu6B/Cda64s3OSNfGwR6Oty0gMzgnpI
ygayr7QcppKewrpuwx6Re7liY5rlanXna1C4t9jdYw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ESPDhrvv6BXab7NjvW9GZy2swPCWYssr+qCHszk0hFhw/XaMcHq2bpUihfb/
nnJbjq5e/s3QL07IW3r8WwL1InqkUoUkyLqs+q829qDajnwz1UhZzROXTOzM
/bEMjfKXbOfovfzJ6L0Yj8HHLz3TyN2oTYbso2ERWHxf5s2OX+s=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lJafp3yAdi4DETFbp0piDhuQNY9r52W0pukOSKPxG56+kj344lMRlNuDvIZk
FRT1V/iltcKHjAzftMNcJ+BkCbnxhy7ziFpm6MmVJ82jIVWT2ysMViDxDtD4
/AKm43RTiMZZu2nB9OIbk4Hqn4873NYF3Cm452ycWBZrZ1SonGQfa2AH6/aY
INK4Jcu3Byuwond8DFuhc29J71kJajtoU3tNp5ldmfxllY4fMzjdeWgIHoB3
Hml0Wa3WvFheKpkgpop6wc9kkkCuGukAHuFe5PcjEyRWIsNxMOuSitXHYL9f
ITCXfSJcpvfICAvx2qY6Bse0/hVq1jQTJbGWZvHfNU5ODUNRnT5IEhh6yzWk
oxdN80A3PGwZZXwZxY5zoaztzYj6xtMfiba2eu4HA3H9A8R/L8GO+hQE60pe
9uBj0PmEfn8hr8uVIMFVBEUWTBdr1BVqLQAYGj+HZ8Q6JK7SDE0TJt26/Qws
iKKx45R7GnoxSxHNaKLKgS5kiB1KwbDK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ngg2Rf2UDAk97oxE0AeAyUIPgwW6ZFHHm+m0bgXYVtozuG/S4w/XLhwKaCBo
PAwZQQM3DbEQ2JxUdcxCHmXAj7SJaqaSU2NusXZRmF9bPbZy/DypwIXFUdow
moUOqRWO8DRe6GEXt8AmzRbRSwaA2XmLTfJOgSG0WZ2WZMKliaw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jRiAlBY+llVR7/wsA2bJW+E++3+M22yGOAcwaPaEFSNjQoKimtdLkK8b2an6
maWTQZaHcexhmkMvuarzmE6by9oQcP53rLZUHQ9tjDWzEpZF0R5QBeYnIzju
YXqxQHlMMXlj7/wTu3Xs24hJW3QLWoEyF2cZLCP9H9jk6rIViug=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4368)
`pragma protect data_block
3SM9+WZhBa+yiiZp1y2f9knbcetVC4pdly+vhkH+5Tpxkcv1IrEt6FqzKbeO
ecjdXPAi2RdVg/E9kodnBxMTWoyZfFv3y2ECHfBd3STuCaBwKRZFuxMOyWF0
VPprxUWJ6fymbXDSqu/iwYQMOeEr91eJ2xbLXNURwVOdqFPnzbLc0Y80RpaW
m40ReHGaJD9kyHbKhzha6u4d23fDGTObPOWDawq9EU35+Kv2GpDCEdBHzP0S
FZxUjz1ZlenkBjhnKGgGEebEIMEVgk09MnGs0QEItB+yf+e8jBUhHMbMh9ax
KZthWuJ3oBmvVfuB9TWCIjbzeF0tCQXpPiEUpk3hlScoeyag3I2P2wXd0mqY
7s0GJEdiO5gTX3iwkeY3i9VHMaCHWyX9sHKakccQc51vKa0Cf0CgoU355AEh
l7Z2nWPlo6nfc1h8/fnoFi2gLnWf6ufi29kPxOu87Ub8QNwJNE6s1P/PufDb
1oDxVqcGp0KPHN/ycsD7KH64F7M0Uaxl8rUm4rI5h/YGgaMMKOw+i9Q0Zi4K
NjXtDAq6zvSXNbfF90+vPvIqd6j6lEujPJsuKkpe408FJsPJLZcQATY4tikP
2xDZgH6ZbInz3b0G93LzTnrinSaLPWHclSazO1WOkdfvK/eo2RXppUoYQ94r
b+6ZWIM3ShXceigC3eCBDY9z5hrGgnQf1NFqk9M3qbPd6p+2jTVK83vShxiu
r4vC4GgjhuPV7bQX5tNl4Ph56IJKapKe8lSUySgVscZfQQR6NGFFw6wh4UaP
giKVzvCeqWHPt2Y5CptBed14RmmkgKlg/PdNX+2KrYEOGvG/4EUdpDFesp6I
fRaHTHTTRAbqRNBoRnLeraU2NPMiQGu8z4Pf4J32lCPYel2UAWNyzYchUnfT
LK77nGxq3Rwakoh4QErlHoc7zHVMjNhrsCFph6/nDuZ2EBXGrxAlI/odit4y
YeOSI1zrFeIW/CTve2fEfOeSOmypzxIma7KvoO/EKRF50nGIBJMxu7sOf673
d235jaeH97PwDpKjiuadUeEhF360OxAox93tfq0KS0vi2FMhV9QZ2JIMdT4v
rpcD2lcogkAsUsW/4hiovQ8NRHYw4RMlI/GtZ3PwAjbm9qFbq84oux9UbS0L
qpcl4ffY9WkXXmv+R1mnvRn1cAhWR56ykTjv3wOy0SSizA86BeGQsC35VxKC
2raHigLhB9RoF7/vwtEp2Yu2jpdkZXe26hVymLE4OutFlbUAdBeiW5PUv2CA
fHvpVoeJWOtYOwU1lE3wj7Md/YFMIKWpbPgEK7b93nX13xOidVqxWFgysH5f
m3H3iQwv3v+YF1Km5MVoKBz1JUKtKSPxR/W92L/zNMX5+TIZj9MIFa80pqai
oRgS0feNy9GLk0VhKdlqFNLmpLyhCYrOQuIFMbtOQ6USFHzyAZ80lTdNI7l/
XTXBq+ub/0aNp3QH9hWTl/aT99diGEzkEFydGF9O/2S5Hnn3/5H0C54ogyve
YsfBvJHurb6nyP3te+YLD+SyVqw138wXL8As9nwF/kMGIJNikdCAI9WCFaPg
EQ8yyHrO4YK3+nO5hEwoadnDO+WhE3fI3/WyInCyQN3G/+u9O7TX+nKldHQO
8x9Zs3cI4qsl+q/IXH6BvwIq84+qK3k804krxe3IOeuCJFJn5VLzPDvzp0rl
72ppH5tzJXSWCS9/fk0zFfoI36r6ishtr/VUCbz+q3Nt5yh9QBittGHh30tD
2w7sUWvahTdXo/JGTQ9ucvAyJkCeznxedxX5BF+D/ut6qgu9aGBjDnAu4mLe
9uWDSF7+g4ee5Pfvo1o/mPnP/ZBhOTZUEdi1GqwjJUTQtqjyR4ZB8CTlzGki
p80zgfEp9k59X1nT07cLJSSBJKHUMIBGgHc0vQ8S1Q2Q01z8Ej/2k+BYlA3a
pEn8s5Spu8gzMabM0+U0iSu/xqMb+w52CX1pyO30wdwcPAtRtCXnEcSzOl6B
fiFILpItnNt96TDAvpsnPqOI9mnvVsIxsoI+/gPChiogLahOtRg8Mqp4zMdD
0s1Mz8jZJs798dbZch9xYoPuDNdi7REzF4AsmGVzZbs04aB4x3Ht83si3K7w
dGYE9fdDJWd5DnBh9XzeAcSOz+0aYie0daPKmDGMXRANZWI16Axtfwry2ZzF
w/TtR28ZqdFqQy9RPFUbrsUwG3mhgstt0bcVlJALatAzNCWFo+atfOJtMd1u
p3J5FJnbU5Z/i6HMbS2ilZA6MBQvBuwKaN4acq3onT7PLQvV5/pIj8aAhXd2
YCKxfslUq+2/XbPn0iwMPk47rAJ1/p7E6nIjIyYadIyUJ4Sp4/y1c08p86rD
9sGZv3KjnLsoA+UVJEiW26Cz4B2cVCOSBm4SzVQeoYjzTPfS0NjZ9pENb/aW
YQvU+Ut/fPB7UPl6IRVDnJe/efKqV9A4930elvkTSe51oyaa1GYDDLrt8K2c
0JGNy6v5ULZCKh6OThXiRi2kNY+LZ1fpbmIFIXY4mtwt6KmZ32TO1K3zSesk
xtxFcrzSUkgyGo2YI+gZgqVEchLSXX6KvwlVlbH8aD1nxWMmfPSkmmMjXU46
3sfSsNbCPm+PcTiRbiZhX8beZXrU3x5DHWHJ4zmOUudFCEq88OlRmlw+yz47
NzrnPR/X6zpeHhumCallOfGkBY5uliIEJtBW92XucUrICzN1tqSM5fTyER0B
NuYFqnFcCjmSE3sksV9cCHViRNLk70wUmkErWe2iqgTIb9frIunMfWDSd13G
v8ocjVeGSEtR67f3r+WxJQqoXALWZai4jhrNVc9DcRT9pMJCNXmgZueGdD9q
qtwN8ZjKXkFgeP7YF/6vUTos/lwks0HXf8mmxf4PH/kH6Vwy98iEf53Rdba0
vlT2bp3R4KL7zY3UajxDuuLudKe+zn5XytaeXDBzlCZ7GlFC7EbhBojlCDQf
QUwYvJjqV1gYQDDV/dh1rmz9lfkns501AbAn91Nno3hHoYHO1eXAq/Jk2gRm
rl13hVvKlfNmLj91tJ9hBzOGHuJyse6X6uUL/7Yhr/fgiRTqd3Gy0aK4/AXe
XQQVeMjLkgs+gNslu84b7nzZFmEeMMWPgMwroF4VqJZI3fV8LcE69UVx2Rj+
cXgIRt73C1kt6ulsK5pF9ur0ny465OoEz1lQavTdzzwVmzl8j8GI3WnCd2vd
L7K0KdEFqjEB9yB58grnPzU4mDoY3IHby2Gn3aqUtzL2SSujV5v1trfJqMwF
CrJRoWD8TrmdSs1MHiN7IcwbXv9ZvdFcjkAVl4pOJtRVpSdZKo0ZH5n8mfua
27B5k5O5XKtpxf1OuB9kWXpfEggDgE9rUFvYI2W1V50rdp16hQd+4X+MbFBe
MW20jh8gas/9p+HfLW8jZyDSG3FpEg19iUFqkmEkONp4glz9XKa4QKcn4m4w
DJV3zWFvJxkq/bYAJ6m30yOC2ZhxpURgA6iRM0nUBND4uzP7g/SMgOmjBvS6
cOffzKtkC+ZludGQGjxSE+EtxNlSzNOd1QgH2IzkhPUQOAQHhQLCCOH+q2/Q
jOIIlmNpy5A1zTgT3f2MgiB1JUpPKE/iuHrNwpLPfK79/gKbcx4VBGvNQQlw
PUNMWYBILkQ+A1FK8Bz74Noq7GZnu61Ne424hH0xud226IFRfNPr6RrSoogV
MiuLKJC9fiQIC6ePXL8ZTqVgaQJjFrsPLsq7GG+/ItdYst+1KwLnXam1V2ZJ
8fsF/Wq5silliK5UNCLZOIyl9o5mTr1IIbkFH15vIswsvxiJNrMYINiO4pMt
SK0pJD6EDI8ms8mG0g8HspFJkxLoMFLsKUt526PqaTk+/N8kugXenzbQfThi
BbiIzuqtijim6BVpUmc/rIU/FHPqLiDHPT1fYg42Q6wgtxSgSxYVnsFoY1UA
M8DnRmrgjZkCh1PxWLmSZiO1DDkB8X8tfddELn/itpevxnVjLM4gPpdGZis6
FcUkbcvIO4QmHiJyXngAULzzldahH6EJnN7wLdkwwLW3puWh3DnGo2SyZLbJ
Z0lzh2ZIYu/bL+E+lHdhdeAE79qhYF9pmvIGgwHcFK5q+i6WRfojE75e4HMq
zu3kRtBrXQhC99KquiDfcahwy/TQZSv4hGDMK81MLBzDyoCpICM986BiGVss
mNwQPcJ4UT7kr31aO9zPR456xVlQRGSFRB9hnuPMO0xPCoFJLk2ACQj+xO1R
8h0bklF1YhJlQnvWF+itg8FguHd7R/mVX6kJFvi9dodksMPV0MP7w1ulUfyV
WTF9VxUBJoNj0VnmSoGy/sl8t6TQpTY/L0nK8ftD3vUNO+/ScLenQZ+VL9Tv
v2UcIguqISM484+/eRzLFnyT4Ixegv5GNxzEaMrcCtKPs1p23lN2qgRHHub9
zCLSUWo+qAraGWHGj+OlrG/RtfNvG09LQ9MjNSTLmdsT1cpcdif91o6wA6r5
DIHFCuhaoC93SOLq2WeHXSNFI0YSgZf1WiPziiqExFbAqYXAYa/rnvemXikO
HWrvLst8pPCN5yDYL4dTCtCz3BAQ8Qt6X6I7RSGdk5TydbZH2xOJrXEgIran
3lXzrgyafgUOLIZUbX7Z7rs2u1HfcpjASqZ4S8PpI59Rj0IfBXHbXg8xnwi8
QpQR6YTfSdBMgsI2YgyUIL1SuBjpfu5lgab2x4xKnAYnjslBGGxdKozfIhDH
RIBPrHhEI6z+MFZHh7o3BSlqC6HLTYSHw74k5HRoU9gXKE33SjpfX9kn0s++
nbTC3P/Nd9pCjeuUCaII7CaQuv+teo2jxqlTYVMofpYtKx0NOAgoeuWmBJt/
qEVrP1GvOYiStMY1nlIgugoXK16L9ne1PFUfIl5kTCkva/zgPgmmsoP2YzKX
ATxFOFKebCEGbZWIFPyzQUiTXg6V/5HSQj8Tdbz66iI8AdRhpEEDUQTqabsI
h3qghw3MVKPLBFCcDiMEfOPiQ1Ryg1bprl/LjmV2SmJXp/g7+fCbZ6+Z6t6G
iSwNHgPZSN+t5eFcsWtJ5O21Y5g8qf5OhFHQAR+H2RrVZ9BkHyP2rRfsa/j4
ppfPOFRI9rarhKWjTNDveebBDXxTE2p+QFi6Wn312nCxX5m1zV+QhyXcDGho
r+6YjIz3y19HJADjlzKDs9lwLSf0UWoqeQ8XN6VM97c4B9c1poHZwBZqgPnl
yxZYvm7xpi+VLHsGrV3QHGECpGXUqlS100LaZe1gzUH56tGcP2LHwX+xqDSe
WuwOxiRdr5aBsAMcFHrWtQPZOvzmwG9AgNMKplgaYxN2e4aulINnvKINEWBE
QKySEoGfh3A0nxFMJhmu1wkp6vPd+Slc9CaHxE4/g09nKrXmOXo3ywlZRJNB
BHj2BnxzTMWD3lldqJggzVG039YJ64DNctTF6JxutQcvEdMD1ZAsuZqKYiHk
rOeOxVR5G/sTVn+2vsi9U7txyD8uTFZ3ZYehphSwBUYz5LuJh+sh8YfbgBMr
mde7e9y2lvIHC6Ffq9a4q71V5+J3/yDgP3z9d0IwM8/Sd2uQrH+yxPqhokWH
Txdac2WaDnF02fxgHIWv/YG5wD38W84v1MM2POZL+nj6DNjfpJsPyUkVgKJZ
p3V5s3bb0ccFzBE7JSzJ9UDf1TQLRmMyy13uBoB9oTyiWthanl1GHAONQ2xo
gS5wPnSxriyCSDIlrEvIyb/3ltOHXKw6mb+CyfVUrdyMTc2r1M6QT9RxEbKe
kGXyz7ZLQsu1xwgfiVWBn7ySKDyv1t9xwMwUKwEZ0XisQx1uCRcyosnfLKGk
X+8m0gLldvs3tcyLsTX2UlueJHbYA4GaBKJLH77r3VubdFLMSEj+vv+g4pcY
8NeF

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "q5w9/+5Kue/STKa5XRRpVGZJHL0ZJeEz5bcA85thYUmp1PIQq+G78CEzW7wlYTXVo+w4BCHd3aSh/18cFjiZbvt4xJJC7ehpF3+ycjY5Nbab8XuVBxV0GtSWyUB3OY5g1z7jhNv9saTklZfq4NIuPRMvUINOi1jN2p9Hk4oe71H1u1YzS2f8oWdLZgHwWW1RhshdKbt99NlJ2sTPdlYrRV4HfVHdWgZ2gEOhvkVbm0tXMLSsnC6Uu+hWYrz9DKbxTcEvqtHaKdx2YxMnSB3BULzXASVcV6u+TgFBry5OsnNEmqsAsLRu15twc1sg81w3B4p4HSEj3ZZrWwBrTO6PQMcIEbb/4ISL5YHK7DtvhiGhN4C0pxoK0qpoa0/853FxKFRj4KeWxTinGarwoar3q1FXvfkq5VZmz1q0GmZuzjLvC7fqqjqKnrj0nfI++OQ9y20R1ZTW35fPIa4ogjUo29ZjoosI1kT+f88PMdxJo9S0DwGz4hNDpiQTKFUe3dNmQdpK8yH1KbeYaBk3KVZHY7GgN3b5BSZf+v/W8iu+dDzt36sK70PNHEysPcTAUPnRZF7zmDo+iQEa/1HzWcKnILdTy1T9hhKTX1n7lwvVdbbzq5WksQQ27n+8qqp3MY5/NvFQbNWKy5cYVQ7IRCT7ZBM1IOUYYqJIpAUH8c4fertS0S1F7fml3CSFDQ76zBgR0OGnDS+5Z6DF8CN6zOGkIjVGI93hw3i2CMCx5lKlYKTKh+tjmf0oH1q3kQuji06dN0f9p7bGWNb1G2LhppDGgbZdgAWIwBZSoHIoZOy7mWc8ADDFpAwLx1vLFWMFOXS7AAWyw35Aj1sb0VrGckruXVctmlGIjYRAXOW/MfL4G6TBDCcUfECs9TMUFBL6wyKVr3Y3GaWEKoDWbQPYMkCxafK5LZYhUblzBEZlsW2gnDIdLypkr64TqwaRdAr62QWeJuYJFoUyaxBoJsXsWBAJuFRC8UB1ce67zGcc8NyrYrNKjkm5ZKXjP3PtiGJZuW3X"
`endif
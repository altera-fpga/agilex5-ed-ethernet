//########################################################################
//# Copyright (C) 2025 Altera Corporation.
//# SPDX-License-Identifier: MIT
//########################################################################

`include "sm_eth_sfp_basic_seq.sv"
`include "sm_eth_sfp_a0_fifo_read_seq.sv"
`include "sm_eth_sfp_a2_fifo_read_seq.sv"
`include "sm_eth_sfp_a0_a2_poll_enable_seq.sv"

//__ACDS_USER_COMMENT__ (C) 2001-2025 Altera Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Altera and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Altera Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Altera
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Altera Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Altera IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Altera and sold
//__ACDS_USER_COMMENT__ by Altera or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Altera products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Altera assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="25.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gar3GdVhuqMAD+ygDleHN+MK52zit41nnAN4+wq8N8Gx7nrwyINpbzY8ar61
OWKVmicCoC4Ihnl3+CxaDCJ88QuBX9T4kLHNTHJMFJ6aa/yUH1hPSUgNAsn/
UVncjob2Hm8aqokm3+snNyAJnngOvE2VmecianVJLdtCaadkYNvhmp61LEB+
VzX0RBDWAglVrEibFjTTu1YCt/5pHC8ZQDcnSIshAoKIOIkDtJYNf0gsOtF6
GyWBl1M6hyGZIMGVUau4q1p/R3hyY6u78jFyXdZDe1GMP449oxKEH16Mg1xe
51C668XClIDtQMAyxIJi9G7x6tQv55LTYdaelXJ+0A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RqznaWQACY0s8qYrbiwl3dVMjdbiVpRwX0U7G06jLJWhUNo180CZPPzRYI4W
j2DKhF6lSq5sK80EEOsdTw7CC4Y9vcIJ0yxpa5K8lpkTVS0mKHSR0Cpx3j2Q
1osMGTUZlQ+K46rq++OggkYp8RbjsSKkGtkOagJMMzc/Z5i9WOMGm9KC92qi
EbCouZVnM2YZQFRXKHPHqun0x+v2pfJVNsyDv+j6RdU3Q43+mKF7++RfaAV7
MqfSzg5s75RmzsM985B2uNrKzz1TY8cwA4JoQ4Eb3ymDv6zxM/h/k/uZawUQ
8AEPeHqzrldgzZytcjeaznoZW2p1iFg8X7qiUtjqdg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oGSWWvl4lqbRD7wl33ARfPAzie2uw9M6KbzSrqv8WWp6HywKeTY4nB1/znbF
ivCtJ+LPxdHP6snJ0qZaVn1Ebf/t0IpHebCJxmV+daQpBWJuhPYdSH0gDwTm
qIiTNOnrcS22i1lE7LEDXtz7A2t5Q/8x0KtUga5+QL8X4FHGHJ+dTS1blpTh
HmCn6urrpZpjz/V5uQ/XjPdzZ8xPUnrUipwOFID8kQ4IkfUNPppW3NHAyGth
hYfvu47YCrjCKO5RIQiz4ULA1jRCRp3V0QdIKlmOQGKqo4wLOrFl1xjbvscD
2LABaUF3R1KwX9Ojb96wlLA8uEOBw4sPj2qErZo0XA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QjWNQDDHUfbZk9f8/A852YU17/JNpAPPw8rySyslekELFGQ/1idf5t3whOTb
5Tng90BcSXEsoPQt0HjdmcYcf4fL5J2xmEuFRNtsRu+N2u9n8+VS0YXg/WfI
PamYveVQDsb3k+7ijlNqTQkHEhbxIHEybAmEsQOL1jfr1H3HbmCYD8L9Jl/u
ouDMYsQ0v8i++APO2+7k1eSy/QkLLEKzfip4+VXOv2rP4x2azRaZU7nXG2en
/J6WBfkwZzEablR9ndrtQoS4TpC0SqlicBDEybkClDzufhdq80z0eGxaF5ct
WY9cuyUIxnL5d/qIJbNB0+EJafs7OgW2B6Wtd6bdNg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qtd9oz6SV0dtIfnFWKwjyforuJ31B5/ozv3z+i7tVNCT+V+edYuOtbogXMHp
57dtcJ4CJCFkBHDABFFDQkmQRITWW0E6+f2X0LW8KlY9VwA+EtZGXfxSYkt3
BbYWKgGoEi514oKMI2Er2IPNf5Bk6KFJuqcALALxL7hnxTQ+9Ws=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bMNsEIZ8l27WSSgSQekPA5bB3/1HZA5qZ8P5J7bssi5fG+qXrlPKsjWSDOHT
Xh4IDgOvk8fbYvI+BUGcOQ4hMd585Oabv7CmK80EReNpFxE1VGaInGlIeGfT
f6qkDC4h+F/ysEqi7TVAc3//Xpd7gdzk/fzD9C+70gFwX5LCkUQpMaA10bbc
2crsikA5TcwBPye8fMvzN7PekYr+EZF7iAdjy5fq67qEodsGtnbLMOt2RPI7
3Jeg0gLw6T5a1NPr2IgxCvON4KpSKxLeDHSSIPsBj5fA2FFcOhPalhps4GZI
qjv0fw7WoSr0+GtVKHbFOcsdgJqaj0r94C4EjorajGR7Y3+tjhLNZXAc0Xiv
ZrSquHqunTb7iYxRa9XEM18IPuU4wDxpL8iOoMj8/SViDmCJP/D+OFZ/KhQG
h3A1jZuLhfumjsdr67V/RH1SwlGOHVKMmOSV7/u4wZ9eCszFSQ4BOkjTHO+7
vtibywy9GDO9OtiWuYPIlzBoOHchBnWh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Kvxcx2F/dIu3+7TD+WysZxot3Wa+4ailRn0DLykf6ntUtV3jMgwiv2xA4nqr
cXDJh0TbJEVCExGho9u9smpGUUXMJsHbyudnfJVYtTqPliQnE1yiPF0mKz48
rYVXfybqTLnLgYm7LPNLcTr09DYGgAv6RF4pK/GMKj++2X+s7ik=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z+fDjTAc+igOGFcX6hNAG6N/ee/e10j9L4amF9g8RZQQDlLHGTA+Qb7cIncD
9KPBYTsxLKnWoNy+4TDWKO9TDLKcxNS6f9bO2Aml0i/GtM9Krq0TXumZ9qRf
W5bfmuCoBwd86PJQpTUM5l0xYrEC8LhCPMMZYuc3YO1A94HJmjk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3888)
`pragma protect data_block
xpW1RuXOc5oYlR8T15thRIOBtzmaBmxDrXUJojjyMF3gZKdLw4qhcg3nA9oh
xOlYKgiyoL9KzdkrKrKpyXZ8YVrCFCS6xn0IHVV9fnGzjZsQ9QwuIGl2bBsf
WlYaT7aTscdj7q6Kh+itZTe2XAHHK/9kGG7YOzCy+BviPcLTX/t016Rcp9D5
M4U4Qmu9k/Zy22ylOftiuojZolmHlvEBSpR0wTtzz4LwrKTrvPXDUUOzHT/x
cFqs17ZlUcN9g5+YRDWRIqi0oUvCocuy7hDilo5ODU50uFKxhb36n8hDjOCd
QSgHHYomM3h9lW/u5Vr/+Hsdj6+3cuMssMf5jOdR4aTFGnJW3d+zb5l2zPCe
tu0A2l86Ze+lUkTvx1kMsKTSua0frKCTexZpuN/wT1po3xByzthllxfNZA+Q
Tw93OHwJ5KQ9Og6arEGotBhNbQo+vNpKTpQYlQ//m73RLp1veraQWEvdBMtN
OJ7J9VmP5nZFKk0BZTyjGigfNBM1+Wnh2yYJyShPzdCXYjSsTLu5pOIJ/XGe
I63VnBjFp4AbvtnSPEgZyT2JZciIXOtajOxBsbuGHNfxaqNeKnmLXEGKHaug
rQYhJnj0H6BytYtMQvSd9czOJAHAm6pED7csIaBo9uNFBRFbNIlurFamGqXK
auQq78Cozbpg+KZyE8ydyVJCuP5xmcPDFtGhhov86eBsUWvRPLfSY3HWgR5R
3iIiH3Zotz9Bd/Lcl2924i7KExoSxOgtYx2ZM8Rf80KRlNsBuag8hry9XwRF
Z2cZsxipfi4TDK2K47VXVk9gc8aPcuy/9eUPLb9JuVRps18uch2K3jH7HpmG
D6fwC0vQwEBO1BiZNjXbUgrOnrwxM0SMMBikav6SBRFN1mnou6Sen4umF9z7
ECdYPoVzPRhzEdi2qZcCRDXc50oNUGXVw3zru0ZxyuNXaY+Wa94n6b5C4dOt
frhzjlDmOuOn8ks1lUyfQmpSmtTZvp5dPezZ8VxTw9OZ0Bw6qJP0CYc8M97q
kGta7Sc/BOCNrk6LSU3dgJffpmsnc57FFyfmw587Sx2dqrULa7aO83LtnnbW
qHHXiLcUAgPVdWH1dTrbdoHTvQ/KAatK6EjyxQfSlp1nwilaJqn5LTaZbdQd
F/zXqHR1zzGB/kc8ISwzaOzQXMj6r7JHgv+pUeCXwb1k3/cjvwUPhEcDILAw
Y0iPSBMUQ6zmcAAlatjLuPn4D4Vk3J5QLDik8fQWc7Ddq4E8PozIVbFjk7Vp
cvzrQNCI1zuIbnTgp+26VfM7GE489KXBdfOUjDs3M3WsJedqoyn8SdUsgnMB
mwt3FhMe3tocVQfX+XqEcI3k1bCwH6eRzJdgiXGcJySwUB9r2lPFGpTfA97S
blJZXy6u1gwZw5gWr/TE6zn8haswMwMpdWiU+PjWt2BISddv/28ysOIzy9Rg
YUAqA77vI9gAbA8MezERLXuQEx8JeX8Ohd2iSXUcIq9QI9FCSfCgMZtmFjsh
6BcHyrdhNW2OxK9lB30sU6U6E1jBlyonZyCcZyDm/yNYJ8xz1bPY4xMAGkVX
4ZYTpt8r6loAoQSvHJP1E54O63lHd9XuMJ9lWSplm3Mh7F4OnpsILCc9LXLN
ua7N18PgUE1J0+BLXlsIOByHBv5Q7Zx1eN/3IXk2RccnTyYHKaqSQnuTsuqc
CNuYq0mw2XW+TP46voMstZJSyd+GfpC5CMuiSrgHq5vyLyhAKErSIHSJWUxP
x2ip40nvbxQ4/SjlbUt9rRY+rfWuqb/ySzXEjRVuB++pqZWG1IOKFJ9atbVB
Q3pkKCkZcFeZ+yBWghPvwKQUWfQrU9uuoquu+T9BR/j9OTleTgSOF5XD+wum
kr4pjqdwuGYCEmLrHPD9D6JiWzq6LuRjK94+sLjFWjKM2kjgD7LtJFURJOJ2
zZODchuu4iusNIevvdltCcM15FppSTWqzh7pZ3nqUGAbPHwshN5h29eKhSz2
4YMHZILUzLgcFu8WMHpI5xAda6FajGrxPZIPG0uqKCn1gCRsSgPwFbqV2KRe
qRgL86ovN/Az/CNBa5fVDWpXfRbIQckW6pCIEW+GDOhB4IChfJZe/bHhenIm
eMv1e/HLgY5hvaKTfMfZ+1hvCToL6N5WRBnedtX3Y0XeVngZOMP6hlJDd7LL
MkFIsFoMfVS5dQGEERanVzYT+TfR28khJGXW6Z5EFcWKXjmoFKMFUM2plChb
l8OJEADvMJd/3dSB0HFaH9YziSFR6cU23OvjIh0bQDLzndWCPdCQkJFtbN+w
w3iyHzV1MrJOO/udy91JE/zsF1x8FXzY21TjY97DrfnTiX301Yx+9IuBFR8Z
bIM9/RzD74fYOWIoxxSvSRjaNzNqQyiYps2nphqnlU0D8m9g8oEm4kj6/7jU
1e76ZPOszeAmwNcCdcyfomMBWRtK2/vwz+iEaQq9NjlrBllP2NQ2k6If/o7q
6t4HmSFUFFNafsrWlPttS1oMi+MLtcpNHUTrXx0ZmeqZMVMHP886e3w/EK5/
u6hMCEa1DfdpTJCnjpldw41prrLCex17KjCoeoF1h6DCFUJg3Rc4KPbeKMTy
YqY8L0hgcwvuQkUcH5HihX9djlT5QsYgtOpt2oHn7kUhbS1z8eqqyIF8rr8F
TJty1H66eiyJ98Qr+7pVBXdCq5yu0spmsOP6PZD4aHM9eoi/Bc4h2GaUzEwV
XZRaPB5tTzlEOr1aj9zJS9J4NFyPNEcKxnHtIAMosjbhmK+2et8a8Y23qCQ5
hghWRuVFF9eTzVIsi1az/Wa8zrgiTz1n1Nq46asrNFp+fjVCATeRsPG5WsMJ
VLUQ1oRCKgImFi6ri9OpbeoRxAuvEiahpRuEOsI8WVWWvHYEAHgoJOi2zB5Y
hM1Pge+49dj2wdPJfTKDptVh3KO3pTwRO2Sbkw7bRgQJHJuHQn/0HNjXLYHY
I+ZlSJducjO61fH5TJNJrLlcThHV3i0uefdZkCzCfl8QcYwGD7xHM9DpkmtN
PjRCHu0V5FljvlFFEI/ngECu+Gkc+GQAaoj3QiEu4b4CQZTkWmwXm1/+dqAc
sczezhOoYCVM64+uAWA9E+VBKAYKBsed2Bits8RBsl+nc9XRGBQq1NXKif0C
oRpB9D/Ko5J8j4M+BL/A9aY9FUVJWQj62vRhHtUUzKzmnxuBHb1N1tLkkwAS
ccvPKJtYe8/29o3MFZ9Eh1YZO8aqqySMIpwpoNOw8jlrQ1h9fG5tjlCpQyIf
FoBw7o3SuVQJZPa8E5iDZhT+IxdVHBJxqNO8/1qRWklJQYjiOsjGeed7oW3y
BAZfTy0aMaKr2hinpu3jJ5bcIGmp/VwArM3C3n9d2fQsZv7OgpT4EMmEUhft
tff6HBJK418jkX2i0L6qrhg/pNIHZ6tPbPPtdg4q4ERjsVb8k3WJ6qCAzE2K
oNaqWTeA7k4sXvIbNL/fNYvCDFW2LPpBxjKSfgAGzmQUoNRs4n7UhqUBx5wE
0zbr+s3pYj+SMn/wZvsdTSBjgTgXOK6Z0M4pcw4/8zVXNpNEYR6wlF3zpLYF
FYL/p1byDFMlDqo4HKs80RT7XBHDuyuaIjhKj5FXA1NoDINZ9usmEJKuGbVe
16s3ucnjN4+8KtZrz8ORGaXSg3uuvHJWr4c5433n3HATO6zeH4Ke5hSv4kW+
ukLgUtgzZwJSCauAt63dApbrQM/ACgJVxzBuJ4xNTEz0g5sWuLP6KDOwJyZ5
q6TE0VdN1WxRiHuFZI+7vCxG4GxUzNC0bFuS6i78yVoTz6GBfoNP4Nd5kW+K
FTeJvrFggk7sEDnvrdUBTUenuCT0o2K0vYKfU4R6/MNvNBcu+v196jANc8+M
a+ZG6tAcyfXTjY24ujM06t4iqG9aVr1OrYJNOBBN1D4AyBm8VmsmaJDhKJ9b
E/I/gqH5Od8hfQKgSHZDEw89ebEHFhOZM1KAPe2Y0T4t0ClprzQRijQ/ZAP2
UazFjpAX1gqvBPJt8FwGIKpo60xhBGkBB4yS70kXE1Xal2SdLoqVqtoKi3Rn
Gjl7rs+8EzpRcPVujPOflFgr3FVoo07igYqRt3nRpgsGZ7rNwmDWgDMmXEES
dLkkqRB5ju1U1I/PMsYpSQk8l0wGAHQ0pZw9RnzAg7pJ52IcGDHcKbaTkyPy
US9eNKlV0J+ytx0oBXAPJCts/67IyeWByCvHtY9MpRwcl56057VYskLvEgQ6
N9vDfVMZbbqqbYQX1L9JUA/6RWd7qHaDczHt1Hg+w5dIG1jbKC9ipAbXi5gW
6IE5TjhQhsRVlaOgTcQbEfwhw/r3JHi1/vMiI/z9WsZgGD5g1nojn+qIaAsN
zYE2rghF0KObAMKGOK+cDVIItEh1rNUqVheQE2NTc3iaF7eIKwU/CHocOwol
uJSAz2K/zPcb/C3wCZfJ4xTsQFS2IqQ51zU89KK/fNcjRjOlX0XVnXC9NaTp
9auJ4u0Zf6rhI7KBVKzOmD0ox3GmOein0SLWrs5SozUQaotNqrHij4u5VsW0
iIceBl9wPt5TK18mF7FAngMClELA8LBVqJ3kzXmr3rzXm4hWkKkOpOdvcv1Z
yog1T+sO6Vr7XFms4Nqixt/9y0jAl3aRXqClYbbFo4kg0wKYDpgoay1QPNZj
wMKvnD3l5dxug6O04J8Xkjqqm7aT+mXxXEkzldQdLM6FZay/I4zWdR5z0nnO
ujA5pJ1MUjl3HkYoMOqDkOFajtODHYBg8YCqcrWUmxtVTPbo97K73Qo7K/bx
A8gchn+488OtRmY4Ffj/6XbSajFuwDE5U4ssQpGpLsoRznBvQYMD6yBGP3fy
yWd+6ICihP/uv5becae/aETjeYH0Jjw5Nb3evedLziep6P/F+h7EdZnnCTKz
t7gi9gfD34KoS2j+A2BqnRnhHGZ3lSdcueVUPWD3LR/IgDGaaOcsguSWzWGi
HqQpO/3cguY9ipCTMwQxsbRI8HzZpEYg509AL29gPFZJQMEfbRmv2L6baw3e
Bkj39E9X9DUF3xVsfoF3ib56PulAVUJdiTYUAaALkTYUeZZB1C8mTMY9Ri8v
60b0CgKXEzBCLGANyLS2aryUrrptpsC4D7VOOTHA68m06NDssdzHz+lUE3w/
/2ocU5lBkdpP24r2ssr90v/k05xOxyIuoHFRMTcKbh2j6b+kCgx9n9HiawjF
r4ZmMBfvQU0yy0BPH5jiM3Hv

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AS4t06cRjueFAROGQPahzFFvh0kY78qjNO6V7UUMbmRsgla7rj/oyqL07jwfU9zrsJ5hFlphHzKrLzsfBNhUNS83MxlHGDt9WdkVGzZG3W6wCh/VsU39+4vADNg7LopPAtnBDl5jhOtj4mkpI7NRCMrjyYgNj2bIAgsiqep8GqYf+ZuygOlmktMpxGeki4rdzEzbu4HWl/nUrWyuEVXwjf3fThMV6ktK/Eu3HgdtrI1toZnXmV619ApuY/NeG8N+sLfjrJduhjzAmXcPgdSgb86Ehy85jmUlGMeQZncftN7K9PQhUZWaBN0CUt9CSTZBE3NzaC/NskTPwXV7jWhOcNgCNafdGHzkrxCfe0qiyCZeAMV8f2yJTdB2NsExRO91K5V1v57e+huLvfKY/JIRQBFFyKItJ8mQ8xCxQVBpAQ4gGIBzFuVwEwi5MJLE+xlxx0kLRhIWvmIygi5LY8oCPdJy1C7kxfTghbX4/EUBRQBf+F8sDgmkjn+sTwRSvtXoy5EE6vVwPxJFCI/2/1jeMSZLuesqPKr8jpQOFzPRkrHtcv8GdzdO226za6qQd6HgD7mZe6jsmqQhg/26PtVdaOEkVW0HOnL/BVBRhKXxRBwHxNwCDHqgXBlPmPaGs/9SWXU4wSIdSncgJDlrq/sdbxnQiXKuQQTSl4UtYEkrdfLbkhZmFL1yqg8wgD50Et1FP2y/JfNcnaeOBXsOJ0rHGHRcRLqJbYwldtjrPqgTLcMFkk9pbqQpfwpq12u2EHuAXDrtQMplWaA0wr8jwcmHKtdhb4F3rPYEYBsh/EBS3P+tgpcVGgrN+41ALz7+df6Xtqq9pLtyOZuqqT2kaUEQjSMwYlEvmpQ/YEzXHwHwAnTUjiM16j7x5pspRKYMDmxF9LTgr6SFDqlylKvxEawJL8xrhlsx4OXKhsqoJSCrXdVueCeoEVQroaJRzeWwPxokyXw9IPlX5Kxs70JTCuO5i6+RNJSgYcM+v5HyzigYDJ+IqDcjgam5016otuoSVGrg"
`endif